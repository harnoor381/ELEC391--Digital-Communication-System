-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
CgiULjNZi1K+YfoH7qUcZI3qegGUmr/Taaf9BbArs9MZmixlEtagdudJrnJ/pPd4DPthVFRL8BS+
3JInfOILoTp04M3WmzPhuX+nmsDgFQtIZYiUVjorqyuh1JdTWcMsBG0DeDQihX+hWWGhNmgGG4GN
2dwdgCR6wQ3yVSAy0QHFamhnjNTcWNJViEa9b8cuK37Hh4fuNCeqeDlstTgg30I/Jw0o7S3GzkeP
bTKcCuEuX6XpbXCZKk2Y1H0/A0VuNsDkH0nQGnIHMLktwy8hVmTJ1lHUcVxaDv0w+85/Q08Wqrh+
tMsggxCFBbB43dPcGBuXEndc4RP8PZ873ZVCFw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 3392)
`protect data_block
o5o2RpdbmuNCT5Hend9FU1RmNDPCaR/d9HUeqGdExQT9eK1AugQgflQYhXKuxzxn0bjsoZ5rlQkm
07DXpm2ZtlkiiwMIEDJ8UYtxCWXmx7Zt9HVHDos73naXx9gBhufKuHHqjmH35/KQrf86IKvieJZJ
TIYNcSn74yNCD+CLqNzT9ujcONyHlECS7pSWHiYoRbbEP9YnPU2Iv3m2486Bbs1ehqhfUzxU10lQ
FARj33fUjtGIualVmIrcKbfqm88qwDIkshtrafCcvfPrFk4b/dEAZPbIFiC27W8acIKnEBDiKHQb
HWXmdNecMg+IBtj44VMCTlHc0bWCu6oz4cJhVvYiK8PKkjd0J1VjPtWJ1tjPPBQmDhU1P/V8Lfjc
k7xDHXCZ2OaZ890JuHrzl6AGOl+0FH71y/4HvcrLMyHmIehhMHirBg4wxkpN8HKxNQkJhVm6Tu/e
DTSXS3KFwPlLMsNE/mnFqzGVCzlwdAZKmm62elzvJDrf0nR+P2dvaZHcPTasHJHYf+e67sYjPEso
jwAr/tnNqcL32c8gCyn2zKAabbqRS/MN0I7Tcs4NQY6q92B0Z4EmZae+oXphIni3nhQQ6AkP6swI
RLQ5acL/O7nPAdQ+RFtdZA4NRHriHkVu/zy8PnHG3vi2Ogw9QJJL2WchK4tGjQZMiVD/6fbBCkc4
13ZcNZjSHI/HS808xdyxw0JAOpyToyvCEt9hZZIFEZAFIzf3Zvdr1bYH42Gtlsx99xWpqNaY+nse
EQOUCkha61xzKSFF4+orqzbLI2X2LDNZ00+N4KoQSZirOnmJDLfPT+qcW5ScBVoWKbXbAjhcRjPk
Cwu3WrGQzgBysVOpnQ1/n6IXE2++3jofQq7bOlN2BArYKSkVrgNpGKkPbySJDVV3/GwWuv9tiR8J
myvEz/K605n0PJzKewSJMd85uNyAkzNjQ9Cwo4LHxoekLRdId+CLV7eAKzrKJ0hM/icsUo4ZbMTc
5HRXX7zek111rPk9tG4bNLU49yh6se0cmd5xiOD6wpkr9nfFqhluAyVbCTcUlt+XOKdk7+CzaI8m
mOtkeCzTbAun4ZP+6ZG1i7BNPdrZEwOP2pem67zJ0E4IFsvCuuZahnnGVLE+pQjm9R7PuRj8G5ZT
RL+WXUcamQhNCDnEU5mxFzwLB4JCVvYiZerFKZU8dgyQN20XW98h64y8E9l8PI6qLQROiC2rk/B2
u+UKXolTqhplHUmMzd5+7SFAw0fIhGJLOP9jHs4CSbq9PVh2oGBEUkRiDaR22jT73lPRTOcedvWN
AvFeZdOnsVjwafnAlPvNwfkS6yu8waYy5q0nn9nA7dtmRAvGb9tWyORGWCFcMAZvaIcg0AZhOK0n
LOTOpDHg6bhJOjZHYnMYu9jlGw4fE/7sXtAi3x/vqCptQcVOvaetFe370yofcRLlybPQ1z3Y+lXt
w23jgt2nJ187wbm03WtHuKMQJSgfvIGcYmf83o6P1YL0GA5gu6Nbc7rK8umoPJ/tWznHyGKEU684
aw5Z4C2NRig036tvJo85mgMLwTs4P3ok70yrSDZYu7RuIha9VLTIfc7GM/BC1TUnm6LxMcWwM2Pv
rqpJwjTlALKYQkQCZC//fw1WidfzXW7YsQPXpTzJol+760E51FmH5vTCKLYmZua1EwLgHpLsagwS
cq7mD/vJ/AKuVJnFfIoAC9280uYnryLX8MiRHe2hyRmWH3SuwBqrtj001kU2lYxHf1spaIeZbr05
2OIWQraPOvFX8pGt2qajO5UqcVDSRoAg56xkxT3+eVFC8l3gWl8UN7etA23mHequHHn+Om1+AtJk
2YNEAgv/1B4M8zei8oZhXC4jhYi3cXcnovBSMK76OU4WjPVFL64YH+Uvf6u+t+jcljjnrHoia7+F
k2GJ+i4B92i0384qpmGSxXLHmoK7Ih3sbb5obRnvcgI3Hxx1RktuQjRcS5p5x2r6fwhGSdjDPlts
qDz3rhOlp7QjLdmJtVDX/5asMIrVzSH+0ptAvzqOGp+basPzlEJzGKxVAuHXr74M/o1+9w+VWC39
KowzwXZ4Y17Dl6xM4siG9PINjCgU9E5eLdWTUnbvIcuStTvYnv3q/kedyIwDHds58KJlzFJcr21A
Rkdwk9n7O3ERhkg7KrQh6DWrnICn3ANgNUlW/w/sZSP4umdLl+N0lQnG3FfrqgnQXf7BheP3wZ/J
BLh+Cs2ucBpcwEQ/wm7OF/xx8bNRtI7jRxifI5egMBQRe3TW6PtCF8ybV58l7FBpI4ETXKp1t8DS
thNM39j/Vo0iJdSn59amTjZPFW3Kf/P5Ewk4PmKSE82bbqErahE+vXI2x6xYh3paUXpumDllOe5j
0J05MpJuFw+TWJEBvi9Py2schhP+XYi/RNcxJz5+fpUW5i9Ss9Itkgwf4VYvvMT+N57jdCvzaE9t
NBNQsUhFZx3AqWQErQhHa2uTgPOQSijlQr922oMV1ePRRwJCD4aYrlD26T2bfkoPpz+SCKuyVm2J
nvvhVrBvGyKK61P9zGsqMYFp711gDYtkpy58wX2oOmsHZSf5qfH1AiO1Rm6RxOz08PaHJ9xUXM3S
AA8qlgHCyS+pqM/oOnx8BiNGNai3USSB3AwncLPhkxxn7Rie6D+nLuRtWgJCy4EnY7kAIXeas4EH
HL6eC0gn/WPp51PI8GHAHo/y2XBM6HjBmrrEpdvVRu+mYOWkM47ypSJNFXKTgg1iM2d/PhTg7hUI
mP7gz3DhzrRCspqy1VB94cMaLlotK3K+a82YjYhapVvJiG1pfEmfbGHCeIVW8IUCgEnHYvwHAK2W
WzyrSCVhsIxdzRbBPK09znZOXcIecG8NwuUqFpo4FsFKrRMFeLiAvROKVpSAcXW6s1egWOFwQY+V
Oob74epY/QDVFQdS7UtgneTWuUs2S8yJiFUuLR0kX/JNDCNgPDKysjjOq5/DShg1IRATPsszJmaN
owN91vVzq5QnSllpy4tQu+JyACITeiV2lMx+Ei2C+tsWeiTFXr5u9cxLTmoKHfjcQQUrKer2M3As
QufrS8sOxVafgmyl8lzu/8x4FiasMhwy6mwkbfi1Ya+GIW2bWIel2AC7gsU+/HeaWUsaCv8PJd/a
oxh86KtLE1mnI6LMDbfDWz7R0lEDAWRnEvdGITdCD9/BYAtZfCGfQhCMtmMYHjKGqBMjLGdT3mFi
KdaxtOmU5Qt0a0ERWds4I22oO6oEb/ka0xN+k38AP56pV4e+pBM59KF76QLYfU0OesDJ/+UnyLtW
ez/2co4c+yzqW3g2IBd7AOrWxdXeYjcLWO9B37iItaUa6bt8NTaQf5e1KzGthUimQh+SX85WUHe+
edsjx1IS5dI7hzanRNlrftjN39jsi30mTEZxzMUmIJY+CsU88QYPZS1VJviJm4fyVkTV/eVoLDsp
P5U/tW0eWSbMXROoB95XrCoRRU6VrYToyIhDOIkAUhQuobY8H0wjuiPrp7Z2Cr2Z7oIyuUvLwhb6
rTH4MSgmcBExa/dVuO5UAfWdDtg/MqXUCjrT+Fnff64iB403xYgD/lmBgoOjPEJ8ykXFRP6prGxf
2wJRZ2KTh5jaJuupCPuhGCfFfloQ5qdOcWk0cXufVTyzziiumwi8Jvreddy0Y8o9hRDsLd1n5kg1
LPki0/YVY7zGOLwWrm/v8SxkNpW8JbhT2wrSd+mjPgtj9Dcg99l7pHqBcwLNKNg2V/upC5CrJm4k
ElGPRx03S3IcDJMn4kDRCPgotfqQ2fDqZz9x7betJE7ShN+qzZ946HRJ6TbhBei6cksVRTc8dZWl
o/wv3yf4SSmjQxlLW1teSGBYIWNO59fNOVZn+/jpCJU6uogT231kFDoUeZq462oS1oOnQCzZRjQB
/OdW17G26J+y1sXtBueaZ3OASXwSBrw3LcEvfNr3hI9wuQyzPTQnYiUzJeOX+ZM0d5SYiWrnuuJ+
xQ9RgGi7/OuYhDCr35D38WCGrw82blZCf7VuCm08CT1JK/RDqobddTNXbiflQgMBwRDqBkCw1l9C
u5x9aX8tX6H9oR6NAg/ShDOdksr2bJNiK2CrTe8dNQV7KosQDSIZBgZcafESy+MIs40m/fmCKqA9
ymgETRp8ZPf+Fg8GhR/qtW5VcwIM2g/k06gD0SzKCYIlShy5742rcbU81QD7Z3AthCb5fPvKzHSb
GRhnDDHZ0TzMImeSgQJrr94BCmwLu6WRDQ9OY1wjshiz25EtrZHMBENTJbsSurHyzX1aH3Xvtm1K
Y41UJrNecbP33Q1ExIEZS2bFqS+fA5DH0wtce27UbKR29BpftwHJwyA+8tECeSyMmzY1Of5etQFH
VDhzD8sqDVO9h2q615fbGzyHMrlJK8P0VwrWH6FvSN6fCBKk+sUtibTsSFapNBbG02lRbkRQtHQ4
xQ+iSAYndBbT8fvW/ulGuE46gnL9zOGZpp33fQJIIVqPhNw0lvmg0/S5cN6MksO3p7ZomZDd9vOT
Fy4tKs3hvqrp8uigS5UCxRMxCnPEBeJVLjpXocc=
`protect end_protected
