��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����,�1	�)��&��(��H����dP7ɨ���:��0����,�6m���Ib� ��JK�yUh^��9���E`���K�
��Q/��V��T�"���-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_d
�t!���N�S��گ/�TNM{�C�5���M��;����L�S�:�{���\p<��)�0W��B�R<Qt��Ԁj,3Ӂ�v��`s�HW��眣�U�Z.͓k����W�z�N��VXi^�p�������LҬ�z���o���1-]�7���+?Kʛ��\������3༇*�螴�J�#H?�9��|��}@|�",%G�Z�s�D�-�1:�p�� I���"סN�]Q���-�!�h�h����>����7�5
�����m3���uqU��$�R#�p��T�M�ɭ�q���v��4p4�;�R���8���<����~.`hJ��Y ��*�n�����<鈞_p�;���X	���/G��>��'�D�7�xy�8C]lr���hJ{�0D��=�?ũ,p9TzFnZ�JC@�-���׼u5x������>��&�j�7�*���h2�Q��Q��wwjR���~��O�ȼ�qꔕ����x���[�)���vn��GV}�����u
���ssg����������	�B�N.�ыV����<�5r�HEY������P�H.[��xh�G����eÖ�SX66�.�0$P�+j��"ޕu ���~�_���j� Ʋ^6cJ�n��M�:ٗ�{o����һ ��;�1�Hp��C��*������l�ܶ�wn�O�e�-��X-s�� HM��4+܆	Un������t���j��\�ײ�.W��t�Mai�vͮT��Y�2�Ȝ🼪�e%B�l9���l�r��������(����b���`a����ݷ�v�*A����4)�9��d۾��ܹ`�S��7�������sꞻ(*�A\����4�.�S\RX���4���FE >bʐZzSWHw����z�)Y]u�@���c�m΅���JC> ����\�P��P��_� E&�f��Gh�/ ê#Ύ<�M2w�q�%���%Re�[B�D���� ��0.����> ��]����p�}KI��w*5;���Q�F������ Y�H�U�<u�@�CP�����C8���zzmWb�N)E���N���UΤ.2m��l�Mi{na�C�>���9 <�J���g���Q1�oϐ�h0��h_��4�f��U��2f?��d���=f~�2����,��6�?K(opl�]
\�q��e��#���2L��~;u#���+����Rڸ@���T��菷���Ǧ�,sK5,�Ĳ��/o"BX�݄\Cc���Z��n�S�]���S ��P�m�ui��mkA���\����j���3�{D��,xj�̡%b\���%H��A���*��A���wK������efl��<���x�/�-9�=RL1��������V`U���G�>���G	4������Frnt�}��G4�2�� ��&7f�Y�jE������.B���1XsW�����78�����y���Ht�"�y�����J��)H^f� 8#�LmB��R[�5�G��eAo䠡 ��W� #�i�\1n�-#���N�+�;�� ��|����д�S9�9ct�R��C�������(c|�@W�`}��d-��c��X8�"M�ݐ�]��-�Ʈ��I[d^U֪<�vv���*���)��k�7�L�����;;PځKɑ�}ܞ,H5lw��%������X�2ǅ���3��[z�)��{�:�Ȉ�*�L�k�wK�LQ�Շh�j�ަ#�4��zpX�yg��͛	�v�����(q�W-�k�n�,M�3�c�m�v���{��u_:e(���G<M�-��իօ�}ֺ]Z5y!�F���9q��h�N�B�r��fM?� ��+M�ʞ�-��/6�1�Yu�I5bo��.���\���Đ��M5}�Q�SO*!��C��<(9.��0�󥪣����Q�t��CSn_쫢;э	Y�EoUH������YG�����ڮ=`��3[��hr(����)!BciS|�\6LOsش�Q�w&��b�!sR��	N�`�)Ԛ�2�5x��Պ��'����ٔ��^�%��A��	h�F��0*����T~�Sgؼ����p� qE�w��a�'Q�Լ+4��@���6F44�1;i:dh!~P�k-N��^π�����r�[����u�D#���6T>��ܹ�B�B����
��M
|�(���Mϔ�is�~�S���#�F�Ohu�[�:�����UG��؞1�#�Ly���U��$Y�.~�)kрQ �\�BGu7IĢ�e*+�k�s��,r�@K��3m'k=HbZ�p1��N��{�1���������F��,r�Q[:�yV��h��4^4i�f33��f{����������M��7R�f+�<+�����"`X��O*�P�����C="@<ǽ�1D��x���t��B�+�	(�)�6:�©sr�ų`v��>0�ÎI,��e&&�M��Y�i��7�H�z�H��q�o����|�#��2T!p��"�Y�����;���tYŲ5O�CF��̀�ȴϗ3˰����"L��j2/�r��90����Y��A��e�k]���'P�}�ǋ!�d'`^P��9���g�Q�|��5[En�:N]-�������]	>Y��_I� ξ��V1C��7��ΣG��1]VP$1A���rP��@��R�(�~�2$�l�(ʁ���/ҷ-�ݺ�ut;� �.ɓ˗m�lD���s-�o�!�����U{�C!�#��d����
����3��� ��n� {ha�q҄�㬭�T��Z��
S��?s�^'ld�ί���U�����UOB�?�C^{�	��+��v�}��C�I��{�ʞ��J�'���C��f�'��{�Y�
Z����������M𣾋����l�`WG�`���`��B��-5�"��l�4�3���jm�r�V�!q�z�`"ًd7
R��Q�
�Y�1� �K�۴��xt>3�m�(�U�\+����@eښk� ����y�:"�e_Mhye?��"�l�ʤЦ�[2��:�x�_)�\t}��b�"���tmE��*Q_rm@�+$��?Wn��:]�WS�}�Ѩ�^p(yTcI�����}�����kE2VAs%L��O�p]��LH�ԻM=�e�U֨�BQqo��~`����c;g1����np&Ij��R�'��p�ȗ[���=��;2��U��~3��Pe������>����q|���W���ׇ B��W��x��͊8s��"�ݻ�����ALO>� �Ҍ��{]�PZS��r ���pM���v��a<�u��'т�+Ov�p��c��wH��7�[y�Yӳ� ̪^'�ǚI�p)�>&~��>uq[����B�l���8�=���Šy`F���n�G>���bx��A������co���=�*����MM������aS�tۉ���Z���<D웇~ l��J��M�߭U'�?�3�FČ^���I�o_�M�k&�����	�����<Mc�ۂ�pL+��S�l!f��D�&hbE���k�cٗNovV%ޡ�?.Ə�x��Y����rJ�2���<>�Jl������}y/�Y�+�. ]_p�/jcڀ�Ъ݁�Z��Dn�z�I�҇���^nށ�c�h��ښ�����°L����)B.����v��(q]!��O�N)sT#���;)&��Rt@.T��I��h�å)��;��"?S��2ko���$�7س��<�nv [-��c���&�VE���ç���OI"�����;�ͣ�aq>2]��1{��i�qp&��R%3|�J��H�T�0I���r�SX��\&�_h�#�(:�p��L�p��Ý�45����@Q����zN���?�a�tZ�a�a��,Ǟ˱��Klv%�ܸZ10�0;��g|j�
�L��<����A�"�'V����_.tv�٧�M�Ne#􀝣='��\b��&��Y���� �#��L*|��O�Cmǰȑĕ,r
�V�W�a?H���Z���Gm��J���8�(����p��w�����8;�!��~���f�>�S���l6j_H���hhh+5 e��	����8w��U@"��8D%Ԕ��bn�����w��~cD�v@FV0Qg�ɴ�(��kJJ�dlta��%[>Lm,ʷ& ��d~B������as�R�F�]���*]F�ST����J�7�#�/��rFb�5kg�c�s��;���*�\h?i���W�k��j41ʡ(8�Wx�N��F����6g˳�W�� 
@�S�}�����>���������\�'G����OY�dq36*����B��+6�Y�P��_K�Ud<mÔ�\6����]R.a�Rz��UPlB�����Q�g��TVn�;��[�� c�y�V��XȈ�@�2#�pP��V�� N�f3��D�d���$��l3������wLis�mX�?ى&� C��f0�o�D�D�I�|�S0(���3j3�%��Q��:4C�CI�0-�>��ds� PaP&d�$}1�h��kW&�k�8�ɢy&�f��mV����o��8����܉}N�^�u��;��&�'�p#��rZ--|v�Ɲ��Q�{b��r����A'���@˭	m��B�����|������wi:ࣔ����ě�U���E�݌F�E�D|��8�ت!dZ��j�aOy�d��;�W!����_�j�J��ц���Ξ*��!��-bi�����q��U��C�?���	s>H��� �8߽�ֲL�����	����☹��ȓ�U��к�"�0�	%�qA��P DI}��Q����\I���Ħ\F��h�c�	�h)��ղ9�Y��Cu���|�$S��J%�bZ)�A�En6n����[~.�����g��R�y�R�˔	N@�OH����ݷ�~���} *jY���V������1i�Sorx�P�[�j��8v�+ʪ�<5>G�Ң��X� �3Ɩ6 ���	_��y�I��k�Y"��	����ؓ_�t�;Ʒ�������؀��(�+t�\!]|�D$��ӻ�����]��������wa�b0���x@�~���Ǟ�8Qcȕ�9o�By��A��EE�؈nX���O�11*���v{���֜}�e)������4�oT�yX��.

�������g�:6���Fx�N�~<"�d�՘w�P��n���ç%�ӎ%`\o�S<�����%������x~p?���Z��~�3��g�p�%������+�vn��9��^E{���c�y�u��]ma������<	���(�&#�l���+%_�} 	WL��<BB8���d��	��o�6ؑ5ޤ�>����:edN���vK��Cdzޔ:	Z����)���5Z�,�냺A��Z^��^�a�4�qW���c��P$�%T|��)U:?R��&�ρ��C���ˬ<�_f6��e�����;����:��X'��e��YG8~���W�O�<k��]I��o����aB*���<k� ��;������zw$�UG0�Ջ���+�@F�a�O���?n���Q��/ё�����>q���������>G=欇��.�V���+�E�` ��;��7��	�`�h��@-����� ����?��7ik�e/�vMq;��x!�."4:�e����x�B�˱�9w���'K��g�l���o�&%Z�>]o5��29]��W���D"�䏴�5$�<�[)Нd?پ1x^�e�̒q�~�q�hjg�w�FM�c��d��D��9k+��t,�ޭ	�;��ȏ�ㇿ%��o`	��2���6��`��{&avNA<Q%�z�g|����o�\i!&�`�T��ݽF0���xz<�f��(^�Nv��Np��J<R����lr�E���VZ�BM�w���-VV�1'���ٝ[H&���<
K��42�E�^��B3N/fy���/������ v-N�(��^�g�����>�mш��O�fk�1���or�K�p:z�,=��RǢ���6�#�Z����4��g�lgބ���P�lb#nW��ԂW���@�\�Q���?�?�9�,�˝�Qwr�]�����n�����@V+��~���8S�k���U1,�4�4B�ŐP%ҥ�Qt.7kf&j��Z3��Z>�(��(D�C�nu]��GOd8��n�C���L�/�.��s$�|��ɒ;)-�4F@#:�K��#������J����3Å�u�[M]��q��3s�].�cƁ%���|JS�At�#hw�UR��ԇ��h+��~!�� ��^�j��� �Sр ���W�V�4�����R�� i#'���k;�H$�&�p������"������٥���I�^C[P!�}RY�+tB��M������.�z࿼d��\o����_�'��Yڵ��Q%I쮧�r5��t?'$ss��/,��%���H� j��!o�f�z4�6�B��?�hn�wM�<�����']�%��>�K�<kn�<��E�4q�.S�.Q���Xy��+(Z�5��p\(M��I��I��lJ�7pzw���D�c��5����}T@̞���C�v�x��S�����I#MF�?Y�0��,���vv�Jm�a�9��h7F�DRR^��בْu�������Q��0ˬ�Ē�c��f�����"7쓍�$��sWo�Y��b�gzC�hsJ^�O�9�Rڥ�iXJ���l.�2�@c����L�	��L �}c���*��r�a����ޛ�°L�-c?��jO���+C� ���G�w������e�?��0��(Ȕ��o�`�q����B՛��>��S��a¡գW��e&�P5��,StW3�Huke�E�L���v����nT�r��FgH�E�W�:�D}��X�g�3��/��F�m�B���������}�fvq�u�I�?j0�w�7c	8�?�D)�����a��A�\qiF�Yx�<Yb��)�ܝ�ݵp��?�̜\2�֧-�˯�L�
�rVGO�(�;��6�#�K���2#>�N�Y�0��I&�\��y�#J�}m�#������N
"|?�(��m'�����>��F"F
}b�4Yq�����{Mz��t��J������<|Xl�]��}�������"��p|�=X�'�e��6����~:��e@�I��	Lٖނ�5�O��Z�/x/�"l��a`�~�� փ�¶�[͇E���t��z��Z=7'��k���uA��WV��_Z�;G�u4�_Z�:Ɣp���Ö��;�����u��Q$�d�b4}�Zڣ�mnK�@����=�����c
Ý�ܘ:b��~�ع�y������8�M��rL�kN>��O�)3\�~��;�h�l%nE}��#}4��u�B~%�p�N��b�GG)~3��߼� ���I��/��l��T�U�,y������z|�M�Z��Y�?�s�� <��V�9ޤ��������#��\r:��e�Q��*�:�Ë���[��/�����ڈ>����w���9��]M���ƌҌ��+y"�N�/�ȟOM���S'l	��ğj�9�e��_�W?���4ؿ�����6�ޱ���E�a>����]4&�Қ-���6p�kZ>;y7y[]�|UZ7�Z;��j����J5��#���	
�B�t���I������L�G�@��Zﮔ��c���Z?�E	
���7�źqD�3�g���IG��`p��Ό�ܶc��j�����9��*�Y(�(
�LS��K\�ׂ��q�Ev�+2L<�������J���ݗ4��jhҋ����w�?4�z��\ 6&��b
��G���x(��&��HIz�:��#��\���2,�H������C��lck%�'���\���>���Ϯt��*zǰL;q�� ��;�囪$pS:�R�Oբ>�F`Y'w�MO[v�}����و���w�1��i��$���9��1��"�$LsU���}�|w���0�B�FF�p�0V.,��Ƕ2FA���n�<��3���2z$<8oH��A�`�fV,���
,�3��U��Zf^΍��W��U��l�8X/�ۮ5&n����^̴��wPʽ�XR7�C���i21
����2�����[��72
�9���O�S뵁	yoWX��*s\G�u�yy0X���([�xN�O%ڟ��ZT��BM�dXO��jX<d�#`᎔�$��Z�J,U��ӫ�<���
Ҿ.�7KsݚJ|��6ZG�V��L�ا��,�R1��+v�e+mX�<.Z�+��m��(H��t�����tOj������k�TS2Ԙ �l)�ߙ ���Y$-6kJ�Fo�V�w#�A�`@� �;`�m����������K@ü�� {��ϡYw��dpd�m'4���y7�S�)aEY�t���#G��P~Ur�$&Ʒ���Ar����[&�;v����+N�SӾ�F�z7z#�M�L� ��lvF�P���*ah,ܽ��<�e�uXB��<V��cS�(�'�6���F�t�V����(����wĀ|=��(�eL��S�E���X�Snwj5P��IGDL������]���+E�
��$ϱb���������9�y\s&27��&�_�Q*���Ag4�
eE�v�)xy�P�S<?@l-7�i��	{�!F>�<xge�5�c��q?-�E��s}�@��Q�TR��u%���$�BR��ѥ)%ic��8B_�����������0��:���Mj����jt�i"�(���A{-�� )�)���p�<�>+ō�C��
]P���"@}6�;϶���M��#�Ky��[EHѕ�$"��b�*���;�W]�����-T-r\%��ʿ����B���^��[��;�M���o��J�mi��'"���3�6����[J�n]�z��{2�T���T�thT���c᪥����Z�]������SS�A5��Һ�3 8iKmK(��\J)�!��<�	�#��Y��躽3*��]��2��	5r�ܨ�N��A��~�:w8��K]W��w�����p��(�	�b%}�]�>۾Sվ���������]���\��mn0���~M�S7S�N�M��I�h���*��'S���Q^�D��SCNs%�8I۞9�"j��lG����2y��2}��sz%���;{tl)+O���;`W�r������:��X�~(!�#��h[�0��4uH��_�1rrV�G->ēZPazT�T�5"��+}����;%�)�w��pbJ�U�O�e� ��9f���r��2�S���)�@uRr�Jf˥��K��M�ϢV�Xs|_�e�0�7��(w	 �?������B��v��/�g���^%���o	�����Hk0���0Yr�@��+lK�n����)�PIy��˴×�ץ�w D�������to�ͯC�������0[�́�
]�lW�^/Q�9��2���nę����/�k��(9)�X�Aw�9m�"	�:�Gj��aQ�]��M�<��^� ���A���ZX�g�bWp�|�B��k�!�2d�>0��)��b�;K�|�<��\����Ma�5'׳%��*
	,c��_%�AW�:�m��e! 	m�a��n��o�,0o��=�`��rx՘�� x���}�G'�}{v�٣q��g�;ۻ\4V���{�2AՏ@(�7��[s�7��L���\32(�P7E��ݖrfc�r���[���¡P.ӛ�D`ٜ�����Z�s�rҁ�0}��/�2�Z@�酹^��Vc�+�+zZ��8��ܨ4<�BS�O�-�����ݙ�����^�S�W�i�ep�W
��^ O�>��֧�ذ���a��rY�Ԫ8а{=�"	�:T�Λ�Q�<�o٠�.|�g��N���f6��V�2"��Ւ����}k�����ޜ�V�s�Ȣ=4��7�Z�'�(�"��Sd9����І4)�`M�#�ks��H7m��b)Iu��0"�&йƾ��/8Sw�]_�9���͋�=ް�4D�|��d��N$�Fv�_���d{�oLy�������C��?o`N��]��l�~���۴����	�����'S��p�nq�6��ai�Fv�,Z��a���p�<����W3���1D�wUl��x5�0Ld(�>~���e�=�?c��q��f���g�mH����Y��`��u'Q�w&��)ߪ�����k"!U*|t�����W���)y���/D���̮�BMxV��옐�}{�= �m��b�;�9�[ V���Pp�`��ek��nwf��Xj#H����n�:�Cs��l>�s���[[MA��Z1��H�N
�u�+���B_��(Dc%*��<k�j��&\�bd��-)�ro�"n�1��*ᓀq���>7��� `�eҝ]}�.9X�y;ȸ>9�q�S�Uo��eq�t#r,�r<�Md�/�+�[�]�O���`��QT5��Rw��êZ���H��D���QY�C��'8@IHl<DѧV�z��|�_��t!��ENk/�;a�����D���Vm�U� ː�V1h4I,5�.Pk�и#�~�$�ZY�
E&֐���H�v�K� A�r&�����C85e_��f�Pэ%�0�0m}t�oM��&��c���f�y���H��\	��o��f��#���&�̶E��3+m�n"�!N�Q0���vp��	c#2�6	�&�� T�K=�`�j���զ���{��p
,�bFE0�;��j��\硦�*��[�=�۸��Z$��P� ݱ��S[¯_�[f�0 c�EI#}�=Rk��͜GS*����p��ʺ�m�!J�- 4��l�jєS}8�0��gW�=�x:4H+������ֻT!���ߍ�_Ӥ��Z����ڞ����TfG(~\�ܵ"����=��%����ԛ�}�8(���'��!9�N~��ʭVi�(��6�<-8V��+��;�LOʶgS�%3�ܶ��G$��Ê(�S�Ḿ����H[=���,|*�Z����H������8�dV���`fN��t��r9��a�Cqsd��h���1����w,�m���V���f;��&a�iݍ�#:��jz�ɚ�����bhyyn�Z,%y����o[�'~��&�{6M��nU�>�+��z���w�A�ԽjW'�m��[��E�GU!W[���-�i�,!��l:� �@@��	���
�E7�,��&�-QZ7�8��f�{����r��Hz0��!B"���v����Z��S�]�;N������|�=��׉��^N�G�l����sU>����������|֒�sE�{MK�i�+(��1�g��qD=�o@r�M�1�[�S�e��n�O^�Չ�kz��3�3[������sn�՞yg1��]�1���Sk�
��OYrp(9���w��kR.c8��cy�Hk�g�	�����������BVd��W��i�s��<k�A�e�e�<�<�hM��0Lu���L׷T�x�X貢�oT��
�Q@x�������q�����hְ-o�63@���?ެx�طɋ������mx�cX#�p��+׶���c�m0	5�
�	Lʜ��s{T� `s4��?���t�E�F5�+S*���}믷�}@�����4ZR?mM_�*�цC����7�4������Z�����|	�{&�-��X:.so~/Z��8G�Ԡߐj��M-��2%F�ס��	t̯�ևI2/��'�mͱ#�JӚ��"^!X�ghmB{���h�ӗ	���_�O���X~��I�h^�I�����H&��UfYH'���t�N#~���j�T�+&L��F_/|�aY���dm���%�ӄ�/^�X��P��5X})Da�O;����;Ae��������]
TH�X� j�߱H���E&|�#B7�0+���#�W�/�_�"Ud�(�@�: @-���CUm��){|�n�䪤 ^��i�4������� ~Y��e��/NE��F���e�����voK��>���V�es�<�m=����zL���cKEl��{W�)^,��ds!�EҮ\ `�Ode�R�?¼{Haƶj��J�S���#��}��H�� c�m�]bF�8!`�rfu��.����N�&E�,�Z�'�,�}��}����n���M�B�{ǳ�M�I�4p�wD��	�E����?������������":�(0�Zܝe^�|�Sn-H��b�E9z0.������JEL]�.��+2�>�ؤ����[84��h����x' ��Zhl���Ʋ/��Fl3U��(�@2�Y�F$���hF�hk���M^䥇���z����g��4��!5L�w�����i�;��0�o�_D�u%#Y7�����G���31j ��Y�0GAE��=���>��4���@t|�������h���� B��]̉+�ءo��@_��!"������U��s6���r�6�!r��1&k��1!�e،��i��ӽ�H0\W�����t1����v����9�j-%v�C�vH���������SI�sBBJ}���)�ew�p���dA��%�$bk��՝��!w�;���}�,eQV�N���Ww����3 �;�c�x �@|�� ���6W�V��:2������O�vK�HP�"m�k������-��F���5����j��V�?τ�]�0�'�����	�ǚr���]��rPE�d(��qWl6�\e��hY���ʜ��+�~]�Ʌ-��߀����u�g����j�%
OuWR����bA9�Z�'����&D��	�/�;��{b[B��]�_��ZZՊ�����Ƀ�C�We�������8�3$���+[5�q��!���� �X��͜d���?�6J��u��P�k_5��3��K���ϒfD*+��*�y�t�+��{��k��5�X����^�Řz,jMT���e��IBR,�H��I����5 Qܒ��>b�N��ͥ��΂h���8���v��$�zr5�\�'����Oj7ީ3�l"���{����n/��DV׫�ףM�|���K�}�ޠ��T���Wc\���+�����	mǟ{��jg/�z��:��X���,�NK���+���x餲���G~���$�c��7L��l���#V��C��qt����fAD��Q��ٺ��ϼ��K[�k�u�?�U���?�*�=�)�A.��3+i�� ��MڢI�Z["�K�ll�׿�̫)0C��d�&�ү:,H�q����$���S��q�)t(�>(M@����
��$��� ��fm]ڄ!���/��L�Xx��H����4��)�|��lP�sz�������w.�vM_�<^��J3g��ͨ��r�-�����f����+���Q�2!�H˃j(Ioc��5�����{�|�}{q������C1��A?�|K��~碎�������<x��ݚp�\��A��RGAD ��7|N%�KJNWu0jf=�}�mܻx5�.���P[T?Bӵ�=-mAlk�����oѭ��@sj�NHS�t�<��mΰ\?Ш-�,$x�z�[1VR�z�@��@��v����񁭝~�\�@n��`����xhT��챼���g3�s�/�������8膱�R���2=� Efٗ���im� �y�/`�Ny���Sk��I�}4/pZ��}�)���Z�"s>�/��B�"���j�(-��h�_W�i���������"��H��i� ,�i��,�2�_����6��H:换Ee��(�H��j\ֿբ���=Gڲ�z�u���lo�C�)]�}jo���{ۦ�C��#~���x\�e��%t�l%n��w��� ��٣9�e�bV��0��ʫ2R��*�ڽ���}P�|��DD3`b!�:��k�����F5tŦ���k��X,_㞋z_��%�o���En����u�{H.0��E"�G�ڦ���,\(���b��5��҄Pd6J�7)�0r��<�Զ�2��T��"p��P߀x�=T�ޟ�,SR3(��ڨ�,����7�X��{κ���Jx2jߛ��j���~�ι���u��8�r�D�>�'qM��������~?�������m�fp�k=��q���E1�Z5�"q� q�a6�{t!�-�x�������ἶp�m� S~L(p�y�ڎ�w�x4N�[\������$Ʋ7�`��yr˦�>]��|��?{ȴ� �ܕ���";
8���x��n�;4����TD�Qc�&���Z?ww�aa��~�|pzW{�=�B+@Kt�y]=�$ç=
��9�M��bw�ȋ�4�R���\�oVR�y�v]�V2�}�#�!?,/���	���2+q��'DE/fa�AG�^ۜ�K����9p�a;OHV���M�g��T{�DLԣ���^�w���tx�;�b%�+@�9�[d��+wi=�9q��M�5ߧj�>Φ����T|���j�8�ծަ"󊂂T���EpK�Qԙv�&�vߺ�Xo��:��C�_��?k*��(��j���5 %���|�Fe���< �ǵn'�M՜�3}�f*$YgQ�Re%X�S�0a���+n1ͲǾ+���ɒ�����o��ݥ��G']ت���@��=�I������;����m��d����`v<>�8=��	8Di?���(b��������J�ש���qyaM�9�%������o�O{�'�:������B~�xg��a;WaB�tSu/�N�-��k��(�-}F��dؿn�#��m��:Τ�$����
Ik��/$�-M�� a�(*�o��d{����5��[@T�v��� �h�0B� �[��X��ꖬ��*T�5�w��1���@�pm���گ�n֯�sh���*ߒ.�s���=�Ii�Q�xH�	_�����G%���7�>q�(�;��� �o��7ާ�Lsg1�СT�Ҳw�뉆M/�Xk�+�F+F^�+���L��d����r>8e���!���!}"����]��u��(O�x�n�_$�Jzԍ�/�Q���_[���p7�]��k���lbU��?�r�D�۬�<�=^��Db^��Z��'��z���>f&��;%�̀�zdN�LtaL�'A.>h��w�����S=��9�y���������mrD�4��F����I�U6D���r���{���3h,�8��ʳ->�,�[��5�z�5͊�qp�E���ƹN\q�҉96N^yrh;�ߺ�@�H�!z���J�]���yP�A.�C�n�fT�^�g���ռ��.j�a=�f�FH��4�`X�J�� P��D����Z�T��}p��ߗH�In�]�d�\��k|���X�1f���a�n��AL�y�M9};��O��ڊ��^���[�N��7�8"qK>���;[����y���/Ǿ
!)�uy���&օ$�/����T�-i������t؋6�����E�}Z.�*��6�\������-��R�/���m�fZ��&���筚l5�� ���'R�f�@�d�F���� ^��ޑ�τ0@ld���6e+�H�r����bߗ�ε���`�X�Y���e'8K��%#|q�@�����t$w�˪?x���)h��O��j��qXp�>O���=od߷Z�@��9� ?���_S/祌K�ѽ3��#�ë���7�yP.GN�2ߟ ^��^|_h��@bW\ًmUۜ����%m�=M�D�Ag��ٚr�R]�OŠrS<w�fi�$��`�e���L����J�&���Q`J� g��g�V�S�!S.����G��{��K��<���b+�=�[�s�JA�����ĵ���`��)"��ȑ���a������c��R�ߛ�&����=Ǵ����A\�RdG��QT+��G i룥���8`k�plT��ɣ��:�����O�.�m�&�����k�����N�M{_=J�ry�F�x�&&K*QI��+7�{�E�n�7##!?�Z�ݠ�7�y�d���&��e�ba���_���[��¦�#
L�c�
���������Yg;rJ��?��CZr��� ���f�:l�K"|�q��a�x����F�z򞈐32]���p�$.���P�P뚡�7[�|��W���aԵ�p����� ~�p��_��j��gvD��U��Nר(!�����b�P$���&e�^��W�t�Q���0�{��Įy茏����|<o���:�xU�.TǛ{+S�v� ����6%��������%�G�c��Ϭ�!Uq^g���0B���7	��kP��ҼT�TբtHұ��R��Qk���+�������N0(��z�js��Nh�8���D��JO�W�VW�B�\[jn��a��5J�+���_��䍚�;w����<��=�z��}-E���,�S^���#`k��hZw0�`@4�H�!�kBE=��c�0D���Eqخ5�%h)�͸�O�+m�s�c�z|79o�g��>،��D��%�G�uOJpӴ������&�fAÓ��������g��5����Z�������8J�6=��6���X�K�;ڴ�9�)�)�$�-���9у4-}�Oc+ ��2�;�G�;�@���+���P�:L\��&�&x\`���j!P��v���p�3Zޢ�F���:�gSF��1��z����+��_\E�|�:[U Uy������I��w'�PRp�꛲"�=en+���v�B�̤��6�T�넣&�w̐Ӹ�q��;�	S��o�]	�&��)є���Ё��� g��1��[�p�n����[�a/���#�c���Y%��#���˜9�kPH�u�� �������+���6
DI>�t �=��w}=�0��$���^~�Z�}�BBJ��s�_i��^��,�1�F����t�c%���w'��f~siz�nj��TRe��@���5	Zg	�{(�5�-ƧeS�bs\u}TQ t�A#8"g+Ψ*���r;0��-ho��x*w:��2w�����0y/�Nv�
)k����c�.<p�ޢܱ��#�h�|x�.Y���l"�����
��&�#�5�	5�a�����;�K��HlAJ�]\��m|e�riA����C/\��+!�x�#-o9������m�N9����	�m�_��C�����	�Τ<�8��,��TYoH�Xo�����d�����*���b8:�	�J��(��^|���rsw*>̊����z��LY/��0��0^�E�i2�����t�*JV\7y
�L�[ʐ��0ڰ��
�y5�,��q��ֆ�l�R��_��<.D�6S�+�^�¬���E�뚣Wű
���{t�J�p���VbG�ѣ�^#��V}bG�W;
?�#^d0�m1>z}W�x��3�RM� ��t&~?�5�f�{�9|��[Y-S��n'i&�$�]/�A�Kk�r=��L���Z���Mc��.�T%b�B��ښ�X�A�]7��q��u�\�t������l�v�r�����Jө��f�J��f%����vW���_yT��[�h��]�y�#��a��JNY��.��&b聛�w�RPy�M��7v!�/<5�Z4ҷ9���<���<���1m��$T�m3fS���t��[��;���WnN4U�%�6�x�����3��i���(}Z�hd�c�HEa4������#%S+ticz�/��fச��T#<넌s����P��p�Bͷ�B�g푯�>/��.��"��)u2�6{�������3y�� ���ҝ9XV����&�0�<�pS���~�y��N�F	�쩃�<�8��a�^�)1��M�3�Aif���$��Y��g��Q��T�K������f��ƈ���b��L�F���$��o������|1�K�	���b#O�}�l'����-Ƕ�(r,�ب��䂸���أ�o;.)m��cQ�f�?=���diL������	�:Fj���N�u�V��H�-��J��͂� R���ˌ.G	B'�N^�u��0��-7_��לK�Ɩ$����Ԯ9����ރă��{�7DV��G�&��	j�԰����+*�m(��M:Ĥ����0a@��%��P@���~�c������m퍶W)k��_�%ݨ��R�[�\oV�՝g����5{�3�k�P�9�z� bR�(x����F�W�k�X��(A��``U������������j��q�Ǟ�Xs�A�m����DP1��M�.��u�[�A���Q��c���jYj$���$X:�	\G��^�%�[>�A��N��O_v�]���(��N�KPcSV��ُ�U!���?!Ee\Z�]!�1�fWi�S�W��a���>�OS��M������d��z���c,+�i�Փ���фI�1m譩�Sd��KN�JE���<�[��^ S� ����w��o����\|��jE�l�����s��Y;�J���7I�p����� IJ�⺂��wJR��Lg�癞1�T��ExݴSTf�p��h��Ua`�%��޾5���b/^�˄N�B�)���]��o~��i����uc�|I����"ʪ�E[E�Q���W2 QJ�ˀi։��$}wf���]@g��&Z`9���y�T�uذ2$��uo/s[�Ǣ�i�W^H��y;ߺbD�<���~�����5��Y���M�i~�,�ۭP�U�=5U��I��'��Iy�Ǯ�yf��)�V zj\�-G��Pvݡϐ���;��<�#�[�<'޽]p�c(�Z�8r١ɉUaʨ�"�O[O�!(��; %�k�� �T>�q�DԼg{+���&�8��@]�	���v�)�K�4���CC���Cnޤ���`$'sX��KF^;�4���̢��yJ�w��	1Wu��C����7�K��	��;2�#�U�5�nI�w�wJ��j����)Ծ�0��,}�RL�I��@ �M��6h�T�v�M~L��u��J�Q�s��Hc�!����
��՚�ڀWY��]-��TR�s�-�c�L�l�D<ɑ���q�q)a18 ��)�m�A���.Ў��%�J�.�ݩR+���ĥ���f�1�����/i�-}��O��m���c�M��+��S����U�өQ&B�ߵP|7��f�(Y�o}U����lɬ�A�|j`��/����:�^�T������U��8m��
���ڛ��)CVζ�/,
��Vҽ4h��ܔq��*��i�E�Z���)�@	\��C�I�_�iw��\ߓ8L$Y?\\�8Ib�l霆݃	�����m�k�� 
qXD�3���+�[�o6��#����� FA���,"��!XG��1�^2���E�g�zaCo�# �5/�4�gzϥK�[�B��b�D���B]�����L�ãn��k߳>�{[���TY�b� }�u���?���KX˷@r�#[�+M/tLPߝ�4ES>�yw����������>	�*G�,Y�)��خ_?{4s���B%��jF�0l��JP8��)�D�K٥Z���Q�5�z��K����e>����_7l��]���؁:+J<��O�ؙ��^��� ���I*t�=�%�f��^;�x��}P�1l$��7���G�+�;���"� ��<�*�+�{�]���brO�Х��!�m��'��v�<G� dB��ۦ"�%��4Z�N�7�Qm�f��G`��5�$����^�eL�����0JFqω&�1#�t9~��0��ׅ}ow}���	$?n\��*2%;��ryR�����G�P6K�_�����ιF}o{E���f�|خX4�Z����a���Ͷ��ڻ�i1?4H�����ڇO����Jc��
H��ɶ����~��͇P:�?(��߀6q��L?'KM!� V3z�&�E�L���/F�n�h���,N� Ⱦ�i!VJ�@�l�$�I��G��en6KdF�U2u3�m�!'4#���`�-~��7,��8`$nJrV���>��؆���G�<4k�^���Mt�#���=��
/�,�R�Ʋ�&V���L�/`��9���̗�P+��=�);�o��:�c؛s
�{Jq&�o�C�~7�:�Sp�C�+b�!�7��W�/0����n.�6�������v-��B(���ߩ�i��GGA��4�����XLؼ?�E�U�-�~0�[p�9��?�Ht�V+�O6Z��jG�P�w��%߇�E��� }������t�{2���Y\��-�=R�J
!ϸt�u�[�*|���Sʣ�S��]ʕ��H��u_am�Q���s�D�7:c9�1�K�s�n.�G֗j�ߢa?� 
2�U�H�n_o���=Ꜿ.
��\�9y��}Eʷ�̈�҂�DB�k'�6�,�H����Z'�Y���zH�5��[�gVW���N�V�/�H�l�nu�F���,���������ѯ8~!9��mv$��ҝ�H��Q60����;<.���lw �`�bH�۬v������ãX��X1�9LK�Ͱ����+ۚ��/�ا"t��� A�3,
�����8��t�pR��C���FZ����9je��?�ˎ��sBې���$��ڳ�:����p�R��K���rb-[��f&A�oy��m��^����Cc8]X��ro�&�����4�b�3���6|t�2d=���,$g����PL#d�hK�����Vܯ6�*�B�쾥i��^\�co��27lu��8�TM��Bf�Y�~u:,�⨟�B<1��r�}<IG��o�5���b��(�'l�es�?<��4����ilX+ ƫt���)������4��ի�Qo+��jE~�>[ԍ�*H:�n��b�$_�k�e ���&w�3. ��;���֤�rF-�
~����y�@z;�Ӓ.
�Ӛt�F������rؼ[��{�Ӏ�0��4ŀ�1i�`���"�q6��s@'7�����͛���Q�<�qO#�.����죍_�qu�MG�>hf�6s��+U���У��R���1\�-��8��2�œ��ǌ�
���F6�h�2���*���]G��&������k�/[{�J=����=�;K3^�ތ/:�5�W��2	�&r���n�]����&㛀��?�;�~��U���n\B��d�ʃ=Q��=bBMC�p�d�nl	����t�)��
�����d����OVҳ	5J$=d�<�WV,�nI�Z�5����-�D��Z���8)M�pL��D�6���H����S��E��}kLѱpx����k���:� Px�~���"���������A혦�Čm$�!i/L�Џ�&��2��Y�'c�eX���3Sh���D4�+Y�+*f�jp�6�r	�o�b%��M��̨(9OW���)���k',�N��;�{�;���\�x�.��*Z42�.g�]��k�ׅ�'�{�JG�,�ֲ�IB̕��W��c�ta��=�nDP�Dji�\�����)ݵ�����x���9��_M'����X$��W_��^B�E59�UQK �[h�st:�x��
��*c��_�WHh��X������p1�tf�����>��kQl`����e��0v���Q�{G�|"�4,.kױ���c����;a&e"�v����۠�6</p�]_��_��{?�a~~�Ɖ�*����5�0e^��Ļ,����u��J�o��f5<6k���'V)f��Շ�"-�NDtR�Ǭ�[��ϭuJ���Fh��E�{�������d��ꄙ�/Gc�nI\܏�rF{t������ɮamw�CG��#��k�{��2vRf=�m2��dCA���/�qw5���G�|���'3!ƞ㋰�I�U��i|ٵ�10TT�`��0s^�$�^:�o���f�H�:�S�.&�=qk�3 ��_ 
=u��%��}�O�ǜ���wx����r�Gn�-4?���j��]�z�K�8Q}i$����u��S�t*�ݞW�2Q��A[ZCxL���p���;N�L��e}qM 
D�og���@~gY\7�C|�.sQ1}F/��D0c/v7}8�_�L].V��3W����ѐ�����6�Q��b[H�/^ u���SZ�@.��B����w�é�9�;�D��0��B�Ѱ� (��q�=@���M�m�+"�?�n�~��n�{�jG�@���'�i�6��7���\��r�}i`�Q�*�#G'mN���m���<�J�N���Z�� +�̷g=��Z|:N��T�a-%��P%<[P����v�y��z�8�d��j[L�"�UArf�^���6�|y�E0X+�^�-\�v��K�h��S��Nf�#l����2�M8p��z�8atK��$mQ��� �~��-vm*�MvޫU�
�@t�)/<|�J�8>QV"k?ث@AE�r�=�D@)���	��R�M�5V�h�Ob�#�3���U �����r���_��2�B�7|*t��7{� a60P�(���+��N�|�Q»�N��wb"������^B<e��o��[,j^y�� i�teВkW�tm�����=!�]�Z���O
��Z�UPe�gbl�^ vH��>ݳ�c+��ܚR�MB�`��-A����S�3��1\gS���q�7��5^�	�ЁY��T��b
�&���P2�X��e�_xSHF U�Ű�Һz�Q¡�ry�$>�<3'Y�I�7���LR+��ad����E1f"G�y�"U.)���}��$!�ݡ�dj��*���;��ʣ��9-��,gK��� �~�Mxލ51�ss���4�2̭�,&R�[>{�}쑡�W�P�n]ޚ�^�iٹ΍�z�$��ݢ2�OѫmvM� ���@��EV	��	'�����c�
�9^���e��1~�Ė��YY�?���${}uv�M�<A�G=�v˂N�4���c�#�1�=���z �lKbA\�[� ����½�d�˒D����-u�='l�U.��t���j��=r�|�� j;�N����.��}�v���W�nqIe�Z���H��8�n;Zc�[���M4�.m�`B� �Z�j �m�S)}P��Ԓn����q���[� ?q�||{?�ŧ�9A�ihCt��)�����6E��}PԞ�����8JUh�^�|wTZ\	\�>�"��@<ep>�ԏ��O����?xW4���G�M�.�����=��E�v�['�-�[Y��V�X%�a9J��	�n��i��%��Q!�pa�gF�����)\��ȉE;��b�ċ�q�[v+7�gE��D;�f_�S2�%/��t�S>�+���K���sbVY"��)f��#�9;*�d)f�M�IaX����d^]>�����zl�LAn&H��.8E�V��2i�CLt�����#��y]�������q�VNo���"+�c��E�����7@ۀ���R�S+;�+\s���]����ހ(�)ԛ��w���������	Jawid��μ��]>6��H����I0;���;j�`'}$���;��b�*�u�g	�P�or�Q��&�P�qw���|KT&9���w�Ά�T�!�V�~ym)��W��7j���'�ga�7�\
�i"ݡi��s��ņ���O"ѫ��YE�}�z�!J��P�����s#�4�p]��Y����L�5υ���e��	$�4�E!�J�?��0�a�M�K���u�ȢI%���`g[fv���|�:7�[��GE�#C��>���rh:���.D��`Υ<0j����@%å�ŵD��V��&�J6��MG�z��`#r=�\�����B��ưS��
��%-����^U�[����V0|dZ�����:�ص��k�iH�^�-�SA���"1�Ҫ+L�X�Wd���%��gw,T����(
�� �G9���i��3�yb6�����3�I1~ZwSU�;+���[�A�纕\�h GlNm8M����<rAx��.�O����� W�[3�
d��ŧ�y�����	d�Bt3�(Ǩ�I�:M�;L������q��i�Ub�i�K���-W�n}djG��rh��?+�$<�W�fs];��u�o���]�t���T2���	M)�"�솙TZ�!�ΐ>ܦo�����}�݀U�b�p�<�=&0,�Vf�C';���*��E�c.8�7�^VY۶S!C�sT��-Z�!��#���`���I��Ў��ZW�Ů�L����&�y�q�l$v�n��2ڟ�B#~�t��NiE�NΚ��`�6�P��'��7����������S�2X$�3�r�8�(�X�	�I'BJ�x7��y7��15k0T����VhL����/�4�41��D�1ޥ/)��lf���z��=��px��U���1� �K��x"�bb���y�&���]_<e�6�x�� �B�y.0b�[�I�-\}�1��EμD��q�/�yi5��F���E n�d��{�E��S����6��#ؓV�c�
�;]��ͽ�pwf&���l Ė��W?`�Pk:7� vH�nK�aeF��a԰�(̸W����K3o�FT,``��<�}�0��E������Ъ�d�~�i
����f?ܑ��;��4��cb�Eܢ����˘G�=h6�>����懽�)2�M�[3��m�P�ӼPM�&`ȕ��8Dt���x5��X�{��iY���W��uu����I���~a}���w[!�JhlU(떗2��4
[��Φ��)x���x�jFpWN��U��#�Yۂ��2^Sv_�ڳ�����d>��
7#�t�KaK+K>�~���)��7�8Y�t��,&��6̠�1�N���0@h��g����v\O��˄������7��ح;9�&�c��"��s$��`���y
kƛo�3�rI��3����*@Iz��%md�������3"'+cZ�g��a�Z������ǎF��>�����X��l����<����z\�!N=����F�|��F(��@����s}�hQpS�h�!'jX{�*]Nj;C����d����wUB�5�p�n�__,�����2�l �,V��2*���J�n��d�lW5e�������Z`�P�,�����s�P'f�m:���/���?�n�MlU��	�4�Y��ՎU_�́��d]ח�wt�=h��	Go?��J�4�hMQ�&P���D=�gE�ի�A��6}i���k�8��jࣁ�����]I҂l��/�|����(sr�����_����ɒ�X�A�'$�ᣎ��Y��^�&�}8c���{�ƴ��rC#f��h�YDH���JO%+���xYcH+�rʞ!(L�A��gv!1.�ML.�]U�2�/��F�)_��i��\˰Rk�Z��jp��)�N<�u��!/�9�h5�F��u������OS��/���gV~���C��k�7�)�2� �7���/T�g����q�#V�[�`ă�
��0��,*���{ʇ���i?��]�7+e���e�]	�1|q@��6�~� �vG��MD��(���A�L�cV��~Zn;�Jp]n�Xm�~*ńcx�g��A_~E.��>z��˞Z���ü$.�� �� �����a��]��p�|�Y���CA�f�=JC�T^��V�U�����*�&��%C�G�r3l��䗙��UI�Ee�L�5$���d��*^��VS���?M)� c>;p-��H~mX�9���8j�֕v{V]a��|uA���t���$�.	J�m�KzQxb���o��~�qt� �"C�evĶ��<�̪D�D��]K� �������Lgo�Д��tke�Pw~1�#�95`��@fg����ĉ��&KAע��z9*�N];�K���1��S�_�]n���5!���ٕ�ƒ�H�g"P:.ee�l��]iT� G�bn���m�d�kP�igr����5_�c���5LY�@�x������c�s�H�uV� x�;��A�Kp�EĄ�8JV�� �^�P�혨6�֒9�i�7}�䂡ąm)��\�K��r-�@��e�!�_Oji�	=�LBw�D<N^���=.G^U2��[��̈����������t|����Q�M�u�:C^%���9�d w����3�ȳ2�)�CE��#U�b��iʅ[�}!�W��&uBW���ߠ�Q��m$'8F%�.�I��.��ų���{�Ko[Έm��N�=�����G�ZIO#U��\�O?Y&��@%o��O�NYI�q/6k���)�!|�m�܆C��1�]i6��aI^NVn_{�c��Q���s�	�V㳠���6���3�`��B�����.�Q�Q]��g�,M�6�l�"Xr�����r�ۣ��'�*(�_�>0�bu�MnuM+�����`ߌ'	
چs�$��%]�J���/���22pR:`Qh֌D�U�X���
;v�e�/�ph��cJZh��\څG�+8YP�Z7�GBS�L_�4����M�;��z00_v�'�Ȓ��H�~�37�����L2ܺ�k�2];k6��TQ�MhjV�c�i��?��Q����^��AZ��< ��.�J�Q7(l~W�=�q3>��C���&�ޔ���4'E6�o!4!�>�(H�Hs�,��T L��.E�� ���Y[��A�ȰR��*����\Hh�1˚����YW��T���RR�g��G��;�F?�R_�[C �����@��'�Z~�aq�6� bI��oa����~�V�a������lxn�_:�.�X�,�b�	�@0�M��f�"A��.�x�J����ݤ�mz���
��<�M���b�wb:�\h!�ԙE�W�4���0�Q8{���٥Đ��c���'�bT�����#</>7  ��7�c#H�l|�[!ۓ���G�t!��H�j.��⬼v����@bo�٬�+���Fp�5��R��-�^u=�3�����md��U�- �)�������1M��R�)~Ў ���GY雊5?�����ae������r���:�Ŕi��P*��y���Y3������Ѷ�VE�pÓ7�C��3��[���3�p�}�����ׇ�( MQfM�����v N�V�ʹ�>�9�$���u}�0�Xq��|$	�L��Y��	�t�$�_��C��DpFz4�N���sC����_�ݗi>E,��aɄj��yܛ����C4��8cJ�����+�q/#��(�aA�|g]l{��W�=�X���>l�1s�ĵW"��L�X�>���1`�z銹����O,��X�(hb�_y�������F�S:��djGx�d��iv%}�D�-�+���'X�z��c�g����Σ��$U�\��G,��U�&
�U�̎6���1���/��l��LnB�nX�/If��Z�}����A��H!��#F:�[^�T�����$|2T ӳ�UU��d����O����,)}ʏ��_5F�'I�w1<�Ƣ��k��̋S�j�LV�0W�l,������%�p�݂R����?�_с5螡@�a�S2�j�|����g��,Po�}n�i�)����)0!YӨ�����v�镱[/��������nɎ!����G�W;�G��=�d���Df,ϐxT�4�E��|$�p��<@w�Hv���o����A2��k�R�?Q�,s��J� ������<&�׈��|�t�w�B�w�-��]�;���pƤ��yx�,{>�]�*�<<Y��@���������(���v]y�&C~�!�>YΠS�Q/3��2�w���g(,�B�4(�GE�I��x�_�N����)��{������c��j�/�`G�)#�թ���g\�����dOW��-�c[K�+{[ �!���/Ҏ�ܛ�x�T�As]����Dv��LG��ulB����I`�%R�z��߯'ǣ��fT(onD�;���:�d-} !�V������cz#�H�`����Fޢ*���a��B�D ���`�-���[�Y]�u��ķ0�t#i�-�Ya�eG�2e�tUy'ʝ�H�a"�GkEؔm��)��6��ɕ21��PypN7<�{�p�~�%���/�ˡ����uzbނ��V�U��n�[;�3����xҀ$���|�ZL�k�����MB�g�W�sz��Iv~��� �a}�)uiNA�ّ� �'��Q@�9�����M��C|�9L�%��� !�e���Ezm��?y�@sq�E9�y>r�k��C�eධ�
{��?���M��p:��A��Y.�����{M��Ey�UʃF�b
��+g���E������@^���a��Y��qn+B����н�9&eP��j�'�§��������0NqP�����ض��d�qN�������=<y����L����s��}e`W˖/&_f����d��L�wK����k�Za��y®f�X�=�iȺ8����l)X�Y�$G,hW�ً��PajYذ�8XM�a�S�����;BuK�9���̹l\-���̂����ېD����с���ǝa됿�f����ǆl��_Ix�@K�|�)�y�&t��g��z���.�Tjg��Þ������0ܷ�|=F��L��f���SU�R�@q�z�~���z�u�2�G��_��!���<��p�'�#T%��)�.I ;���B<�:��M��йI����*���Β��8��Uw�2�ky��:<�h!P�̕~���̔z$�5�Uo���HD�^�@L�_ʆ�ۋr�߱b�[�6�W��2 4��p&�>���GK�!i!�"�����-�܎B7��x�}�j�Cԫ|h:��\j@5#�;9�Ց���Ql5n�1�I������p�TdIǠH*���4��X�5f6��z
r�0L���g�ci��e��J0����|eS&�05	�5��pd��f8ԓ��%����q��Q���#�\Մ�6m�%�n2���
Eղe=��$�_z����9L�nU�]Ja!�����L�Y���e:I	|r7��L����z00����{y����wt���}f*TM��4f�ML�����t���W��l������Сe������v���=4�[�Ŵ�������f�'/1�iY�c�;#j���Py4w��O�B{z��K\��.��!폙X5M1��̗�ԇ�28�3�"��/�g��"���]��â�Cڵ�6S4��k4n��9�+�D������-��J������x_��)>��˒%��h�y�Zw##aui��G��h�Hř[Q���'�XIS��.���x�[Jr|����G��!�[�m�����|q��9�;�����-"���K;hzt�
��'H�{��:����!>1q>��\&��ۗ³x��X嶂$(��i��(j��h[��{��79�~R-�FZ	54;��$;�%��c20�P���E �Ŀ�>�ߟ��+�Whⴋ�͉7�|-��T�e �.�� ����e�ƹ۹�@����(�p���??m{����3m/� �:�1A���D����C ��������cF����R�]|(�+$�F������N��U�Kg:�+���% 7�NB� ��Z��?0-.�&��9����>��s_�L��������[ǣ�1�(J髠C]�+�@�N�@����F�ه)��H�9S�b�i������W|�s��[�YX�j��	�Gq�E:�i[�޸��:T� �.li�����/�ynYG�I���+�2���lqw�g_E��|����˝_���S}�}�{;L������ҎC�$' ��V=�٘%�^I�\7����;i�',�e��ѻX�
�7��:���kގ)�D�����%�K^S�~d�{��[��ƺҐԉ���I�16ΠM�,;Et����3[^_ݚ0�����;!.!�r��6J�s�x4�4ZR�Ah!���Aap��*��E"��	O;z���z"K6X�l���R�q�߀i�O/�0-��D��ҏ��k��(�=���,ɾ�[�G� Lj,7�ͯg�WڣI�����G��BlW�h�)�ku_���8�`��vQ-�ǒ�`1�����ch��*���IDEdK�PbG��(���~m�ڞ��XLE����}<jٌx>S��ʎx~�ȏ�+�Ҹ����[]C�н�-��M@VVBf:��K���(���b�y#���Q^#�C�A���/��eu���?��1E��2�`�(K ��[��1DM��4g�kā=��UT��ADh�YP��.@Rn�t����E�})�V���S�L�����!�����H�����}�Z;]v��fcr4�"��^�SeC(�(��d�WD_��"3��H<����?&W��DvXY+�(xO�������M�7�N����[�@Ҿ<40X��e�ɶ^����S�g;1=s�����3FD�Mrǐ���Y�m��$7䲶N'��t�����W�rP 797� �W��7��82ʵ�Z���Y�[^�4c�Y,��k��luPY@"��+/(��󷷴{�;��������K�1L���+�I1cf�����%>�
!C3ܚl�pߠ����˱��Ιa�V�B'��l��q�@�8�&�Ɋb|�a�~���pkWu/�ˈO}�6���!���}���|٩�iH������ c��/�x��j�%x��A-Nx���^yRA�[��a�6��Y��x�����ǯd�ݰer^�/�UA��9#�m=e��ΐq�ܵu�i�� Z�b�cG ��� /�.��o$�K<���hTg��[?�p�e�
V���Fr��G!��,�4�e*pqc�B�Yi��hW�������#�!���:��ʷ�x�@$Ԇ��:�Oc��xA;JM���8p�$��y����܌����Y2�D��#_��l��|#ApCū���ѻ/u�YN��y5�s������9�N�������UtC��;���~�;�v�^�HfF���|��b��x��w�D$�t�qO�/Y�F(S�����4L��ϣ�T]5��)�Y��p	������?p�0�޳.�'��B�T0v(y��a�{G5�1�O�W"QƅI��g����ի(�����*0�~n����S���u���.��GB����&sIg���"����jY�^��%^�Bo��P46��,����jy8,Ak�4,��E���n��%�1b]�ƌʮ ��:t���Ji�������HЭ��8h�6o L+�Vh��Aݶ;�hB��E��;�dQ�*\�;z�W;aw�gA{w�}���j�SQ�Q�n �s�]U�)Ҽ�"M��:VYي�}V55��P�s�����\����JJ�c;r��SO\�d�K"V������SY��ǫ�H��r!��h_�,�@M7���g�J�>�ӱ�`�6��g����)�e�_2����3J�wt���C�خWX���W�E�����l �L&��	x΃�@q�=*��ғq�����!��+�gM�\��y�j��K�d_(�п)K���+&fꔠ�+�ʲh�^�C>�L*y7��-�mΣ����d@����{֚��z2=#%�	ZWAG�>��_��g[�
�!���Qxi1�y|��\խ(�w�+Y��bJ�BT%�c��<~���߻ ��ZU��?{��� °�$u��0-lŨ��|��j�dg�W��3uY6��(���뙾�^�/cTz��k�,K�}�Jn-�l���5��G-���,�~�+�߲jR�H��pϮ�+<�3Ċ��-�.6[�#�]B!B!$Kcl�[갱�T�0��P�P���,�*5}%c�4�Bg*�$�U#0�T��`R�j4�,���6���'��х��r�V/Peʊ#r)K�l��{�Q����`��ˉ��j�,|�x\�K�Ӈ;<���s�|�p�2�(�b�3�t��H�Fa������`�r�ɤ��O���#���";sM��n)L�'K��"��F������ݳ�L\�i���0�Fo=��z�'��6����yx^R�g��;5�b	/.�drHS֝0Q��W�	�8��z� ][�LQ�;�<[�������ታ=%�jBzB.��?պ6�9�߷$D5��$� ��ǫ��RGK�0�I���9Ⱥ'H�,�|�l� w[���xb[e��l�����P�X[>k�IOU����
�S�&�&T��x��Yq��b�}���$�x�r{o�s��G��'G�୩�:ڀG��j�k�&cJM6�'��OڪKJ%%g��H2�Dw�;&�ە?�F�8���)X�ÿ�L͠���I���_���-h ξ�6e���Z
��W3TՉ�($}YY�7�q[#�T ��҃����;�̇�&��q��K.����T})mCo������Ɔc�B�q{����`���� �V�\��7��ǜu���#
jW@��z��BY�	�q�zR�(��P�>D�{�����5�%)�{��ˍ�}P�~I�ޕ�<�Oh��?�i��%Gobk��Uw{@ÙW�P���P��;����7mUڳr��H�M��鸲�e@\ ]�a��#u�oF{���Ed1@���>�QP�YjBV��
Ǥ��̈́���T�����g�4w��Q�ښ�<��v��ܜh�s�Lm��[sF��D��r���N��Y
��_��0�έS�Ӛ�C]���u���%�'�[pt_��C�i!ja� _
�%q�95����0��{`y�U�����Y�w�*L�4�j��Y�d!�w!T�9hh���4������3cNsr�^
��pr'Ҫ��±��E���o�;�P��&;,,�K�S����i�\Ɖ�ϛ��bGs;�#���9oH�֓�j��G��5�2��N��v�@iv�ژ�Q�k�������#��])����.g�
N���W��3W�~]��ic�!6+��J;������&4C[��\��B�o�w��ePX��i���l������K4�ǎ���X���:A;�'��x�*�Vo'
�4�`87�"9m�j �O���z��?CW�]L�p�(s�d\RE�+���
9�7b�H���"+��
,REꇛ<�y���VI7���ιCi����j7�V�Y˟�́��pÕL��q�C�G������&�_�7��?ѐk�M����g�'^K�~��<��0ڱ���܎��"MUθ}1Q�ŷ�[�I�tձ�cgЖ���R@����e�zB��<���󊂼����iC�s��&�<��3d����^\��8���k>55�2=�F }*�yݽ��즍)^(�� 2a���:m5�Y'�1��OD{��G�Z!�)|�`�z���ow9~0�*��������"���3�&�Dխ�1�P�����,Ď���N\��V�@k�Q$���Kԩ�B[k4�lS����5��T���<�������l�qp7z�ri�9����
�\9
9F�PcǤ	��D�g$Ɲ��OT7�2�;xĒ��b}��/���:��-#Z�������T�4#��U�ݼg'+�Ř4�P�!2���ļ���q�]ױH��^�+#��6@�ZtU���(M��|3��i%"1��O��]|����s���%��d�ü��/g�@_�2���{l߇�?�/CX@�6������4��X�a�g�H u�;I�fe�\6��RG$�nk�G�a�Q�d�aNW�29a�%����]��	mi:�7G�\��HZ���?v��W?4Zh����7�W�fn�Q_����;t���YI ����~<�jcKݰt���~�CC?I��C�[���E��?���~BԬ���f�9Bɭ��k�0)���5���;
��1��C����%������в���=�hRz&��JnZ��x��%���畂q�K7��?y��T
WP,{����F��iY3CBr?�����̭p����`Qk2�� K��P���?�tFZ=�)��h��?)L�8ˍ'���5�]�'� �np��M���aKٍ_&�z|ƕ�#ʫU��52��>��5؉�������m�p@c1ۃ����V�%߰l�lXT��/K'��kׄ�>+\Ԙ�>Chh��k��!oi�ʵ�@[[��R:�O��er�b�Ɛ��.d�~/��z:��q�_���`�<��f����%���SK̈�hS��zxH��l�GO���s?�2�3u8��B✃��%�#oeA~\�
/)�L��{�G�s�ެ���a6�v���k�ɿ?�MK�� �����jM�+�d�-���E�\PNs 2��`<e@���8���@�k  ����k�[Kp�H���j�>t�z�~���u[ap/pI]1���V���K�+dH��#c�cU9��/6�n�F�؉��	A����J�����9��:K��������#I�F����$4�j�Nx�{Ҕ�d5�H�|
�%{r��j"��65X�!=m��$b��dy��`��3�N�+	�읕�E�ҹ����W]k)�z�[�憂�N�鰉]�U��8	�F�gt7[���>�6+���&3E@Hø�U8v(wҿ�[�k������@z�Wg#����b���ˤ�`;��n��`�0�h�Z?O�C'��t��eS��D��nt�j��.��PA����PSob���h����G6�� �$տ�BJ�=Vg{L�XS!Xn�;EHK��bS��>�h�/c�"E]P�ز�������?sA�U���ȡr1	���kؑ2 K�0��������V�w��OE��F�C,�uC.gB��6Y�4�|^@*{���5`�u����&~a�0�Mxwl�{!��ǘHe(��ي'%��:d_3@����ಧK2������+�(HF��Y�P�J��BF��N&��E��}��2�!?�9������&ڽ=y7Q��r��d�gA�ܶ{Gw3z�`c�'�9AC��;<u�����6�� #�J�/W���2"�][ ���h̽?�	�F�eUSv����4:�MI�~?KU��������q�5�:.��LX�L���n��� ���'c�[���]r�d��#�n�t�YB,E_R<X�䖬;�慭3�Rv�r{(�C!�fk/c �7����OU_ ��I�]�뛱t����zf݌�#��RQ��p��(t�9����X+�)�b%�0Cu�X�:%���qMg��%�]t�Yxܦ�D�B�("ڲ��]����f��z���kõ}���A^�O�*�#lYZ\,�,���Il�4R0j�5D�4�L��������!�y�`�Uo�:���wP�6� �Ƹ��}^?��Ƅf ����9K�KSn���������F���#D��GmH�g�+�փ�����C��\0k�1&f
�U%v�����8OB��7�g=&�	�$�2���ih���kH�b�Xq�*l�Sg=E��X=�rpsK�Sx!3%�P���+���,ڍ^��SpE��[�{x�W��#|k*��_�:N��
3��A����Y<��7�.zmx	�d��h�c�,$�1ϳō�50o� �P�*�B�At?a��9�ۄ3�y�kcԄg�j
����!����|"����ʺc��kj���٤f��,d��u�m<1t�;W��e�Q���-Gf�k�^�Z ����^����h�ơ+�Hܻ�}Kީ(����ު�1�����K*�Wz�>@��c� '�t��9���BFOY��O�Sﭿ�^i��
�(6ᑺalmtq@�(ѡjRR��[�����t�X��Շs���G�sR�َ�&�E��F���~=|��ˠ%1b����Y�v>	�k� sPw�➲3=�I�Ƴ��YwE[3�Ѕ��_w�����c*�袌%�x���Xp�GZ�ȋ�hr���a7��8�HXe�����C�����8{F�2Ø�Sࡺ��ę��ck#^�����:��C%��w<�9k�P�}7'�_�o��WT��xJ���	ߩ�۞j>LR>j{�%%Ę�e�#�|6Վ��k9J�;\S�j_ 1���yLĀи�Mi$���$@����-�G���w��\�J=:���R�������V(�(��3�zog� T�K��Nو/ ����:����P�X�9{W$�,&�<73N�;�o�'�M���_6jГ�X��{�����	��8������t<�䞂�9�t��w#�'m��bN��{lK�zm�͑����0~�wd��0vI7������A�:B i��zw����/8�s��鷹�F�1���R).�ɰ2A���FR�Ͱ����y�ri�{�Cw6���#OghV\�,v����A+^��ڔ�mD5e��d��cǶq�|��3:�zR97X	���̥�PDWU��*!E����>�ˍ���􍎂F���h7_t��'�H�����(*�Tΐ]]��/�mN�t�4���nF�m3Tv����,��q����|[J��H���}��F���F1Lԧ�ߴ���C�ʵmU�>�P�k���۬��'L3���Ť 1_vI�'ߞ��
����R��1r��^h��gl��ހ���!
�eI�����q��]`w8S]\�bE-��E
hr�Ѽ e���ge��3O;��ʛW'�������N��бtR~��/@�,����B�Ͻ�z<�\P���Y=%/����B]0݂�(�+Z���J���0��h���[���fh���߾8b���9`B$*_��6 �yu��J>�����¸KFV��;/�>��g o,[|�j�����AZ��-�\��l�3�ﺼ1S�(h0��.�������C����S��
�*���{�4��#�OSGX~�
<�g�ވ��g�(:�޲F��тI��Qٱ�5��9J�z��LFiͧ�<٭}��D�Y*2��y�xB>2��!�#G ;e��(a4��gQ�ɴJ��	:���gVp�|�A>�3�R~R-�"�05�2��43�oF�w+��݇?���Nīq�8ha��y�x���T�#���s)�uja�l����Z�����{�����AY�q�a�4�x�-I	��O\�&<щJ+�8�)����I�����p/��T<������Q�u|�Mt��2xU����;hg���*��F? _��W�G~��g�����!`G����q�E4�=�;�4%�7t��`�6 ���3�E�� Y%�.�N/Ѵ�O���,T�^ʬ��LJq��3NR&]���Ψ������ԩ����z��:�g��+Է8u��