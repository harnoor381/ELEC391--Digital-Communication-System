-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
mVUkmVfzb1tkkDzbV3S9ZuciFeBaKf7adMTaHHXJ5Q55M+PyFSH22sbSQ3VZ3UU/eyXn+wBQXRzQ
bnhNTZkfZUElb92zsHqVf/XF5yOUm9oj8+VSYVKVPgkCrF20vS2PXThMjYjw+b1VRlbbnoNgTNUs
wCh7ByIq0GeRzxtYZXvjON0MPrcayf0BsnD5UnE4QHi6V0SxKPEAnP/TjZPMjmH0yUTqWIuhztn/
wH3UojehZSoflGAwksqICBksN7QhOU0/KrYm7MT19BuBpY+eXxWRsVb5xG4juA5A62gX70fVflrI
T5ZewmwGQMBrFpC9wWcVwWH+ysnT5tQIOBjHuQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 91392)
`protect data_block
LTufepZ0S6ltt+VsDg2XKFTk6AugxWETo3TWxwepFKzMdclG+GxAU3oLSOumc+EUktZapbwXqjOL
Uwrkgn3Def8IC/tB05vpQqFYpxEDtg0CGUcPv2G+uAwDKSQRXBaIBE+8gIBWz9gM5G+lJXFIrnN7
2qDmDuGJoMQjXLpQl1+KEOZXhPV3DetD45jd+ycIHrhSmP/S/nhD6K7mXhocFb9quyAJKlsM8pau
6EEMURfc1UURjHenEN7YPR134CrMVipo+1qdjCUVSsCMlvcqg1xf7RFcQIrTu+B3yH2aBrzcNLOR
YvO7bEq4nDdazEpLSeC/T9rRVJhlY4vjEjh19+sCnr1I7ig7W75p4iziYEaM3dkknDO7+sRSnkBF
ureiMeVEHVLrFrL2oZND/bex5S7e0ZlU0oEQK6aIEJi7Hniwkutp9tahj8bxq4LuSkAx2bEs4TLN
/z3uxvofu91/agq+5FM/g4na9GWBYV/odUJFeCPrj4d8TJM8kSWPbgdfp/ZZ2NDbI+7Uvyht9LHX
vXSG6LX1t1cAV6302QOPleptY4ys/ffRsktNJGwIpK1Pprf8Ya9x88IcBRsJrI2YOWwmIlj3UJyH
wngLGIAVUULg+TBJ25skM1KmdxAky8CWhVciMsrMi+YVA+mzOHnnsWDntvXE/ycdYWvKlrRAuFI9
vORYHnAVLloC2/raZelp830iTxtbcYGoUdmDlTAxqzF2Y5wwtNzKB+8j1Xn7xg4rzr/rn1XoDm8z
ep4o5XoyYpmkkH5Md9xoxUsDVAuctzX7mlYif6XBPEowFFS6dkoktNi8lWa6TgBHhBGdCX8TfUz6
HHiZrh4xEQVkKKD7G1XJhrKcqroHY0SDelkLlxt8e4UjNuonsgBrukWM478t5JziGLhWPNItj9No
dkj9esKjNuxg92uq6sIENtUUnD23X9BLZApBuu3SdQh0FMRQxqRNwnRUi0h+jVzGg2ea2pFK7ypw
NO+mWx30MGTH24L+9Usj+uBUCNf0fTodGz7GtZn4sE+0jiE/LOMDsKiAiK1SnIgSF8T9bT2CWBw8
psKNugIaIVjFGjVlbnsl5FXdyQZW9G61pLqnktyU/an1V5wN1QoLYuq52gF7QC9Lx7MHAjY29H/D
fJV3mwGo/GYTBjDQgi/k2NbbQke6PX/46rw+5heGPLNvoRq+CyDBHIUEF0TSu5OwhYvR0wK7TIwM
SEPTkJTK4rlhhJyYBC5XTsQIoGd4GCl9QSOy3CDRTGg5Ans5fbKKntrvfM14gdRik+a3jR3VtFLP
SzTTkc+GrTUKNKTJUiC6dOSWm1FCRtvbmY2b4BAWMIqMoRJ5EmFKLC3qMXLClAzYNWoIXQcL2laV
CNm5iX4DS3phj64Hq5Qlg9lM++9EOGhITaCsWOHVq7i4C44NIM1hV9DjOuM2wYaAEJ5IvCkLqHxJ
vjvMLsdvXs3VuSUKP1RnGeSt3mS7X6EYO7v8p9EM9s9vpW9y24H3B+0KuEmT9gdJtdU4net1uuXg
Ho/kJHpKk3iQZVgLEEWodX6oNACf7Svl6ZVpDV7PXcQ1x7W+3J0yOU4rtngTbQQhLHRMTgS6UJ6k
8j/Rwj6ziOw5gLTTXMPkvMvD0xMe3vePpn1L0qstNu4SJSRFHNqk+LGkFwZroSrjhS6RiNkxDXgc
LZxycGhX3xqF+orm6dLHDaiZc48fnllTSueDOs1V+lftnsIGxwNta9KzhUaT4HS1w8iwvRw0PhwT
uOECrM7oE9xkQciLujwSRBI/EUyNuLCNz1rOWLFf3OpVl4V4KhIJEkmm2FmnalptS7pjWOIJpwc4
tmQi0M8F3pqZeaugiEtE00PUGtL88Wp73ayQ+yBCpzxxhn25HNYVQRxU09dTzYj/T04ghUzVrbDb
H1+i9fOljIXqCGnTuqIhpRLc/tn9QjTdf/wp4Oc/NBF8sl8NPBTXi3oYjSQMlKzXn7dpGUvrhdM6
H2xGT2gPMG8j++Cq2niWTwQckw1V40l4+KWhiBIKiZZEtz8mj8P4xC8SGSudw2MIx9gUUKCWoOgt
UEF22cQZtcP9e+A5Jy0fRvM7XBAPrlOjlw/6zzPYLJxXJxR21sVKECZIucXTF9+xRqop4WwsAgJq
ZiBh6uKohIkV0eW3nwr6lsc9ZC1A94FbNjv+DpmTtBwhhsbaliU/08lwJL9fHWyPYrtUvriDh0Pa
nkRo/zvfYseb4klVreXt2IOYhgwBFGQqNmNNzXxKWzimHK6zT2fO0w86fNrtn3aJnjvEHh07OYQ4
f2b17nHA77kwZYQ9E/LUsX/XNjRj1kRqZ7GqRcs3Fwpm3B7w1uKnW9TVS5y4mAOIDxpMkOWXPhJ4
/uC+GuplarRG31RR60tWYYzW2/vQTmXIIhxVw8RM4nOCLzwNvCCP7o5O/eq+bLENE7gLkuNPs84R
uSv0Y8qH4HsklaR1eLw48mFrJHgFtEDWZ/qPkyORpkHTnhEMZnWvsX9INGxjraCR7z2u56daLkoQ
vnh4oDWI6FhRvIKxv3VLVYctD0nXYw8Zsq/Gt/WUIcufpGi81PaZg/HVwRhKX86iPR+ykfCmINoy
BFEeQ33Wc8vl6VXrlA4Bv20Ckdyycj5qnWCV9Bklza5Y6SF3Su+KwL4bIuA5cPkTDKYlcWNldaDS
zFLa8+aGd8xzpjnor9FaXFYB/y7za8vLDpwEcqjnXlUxYVkjtCEDOkeheAZY6JVkwkfDqESQG70j
rBqM0nCJWqtx7s/CkGKZE5npO/MWBFb52QCaO9jKR0K2U9yLu/c+0o7bJR+wcwQQEGbhMU57l/jM
QlItTbuHnBrhUYVNJ6J8+Bc4jA8o5EMoEzlwRWuxZr+OnRDzyDzE87kodQTwrd20Rg6LKUXKSa3R
SKRT+2Pb08fs3zdw5YMdPk4aNSlPNXcz8eHXmYKqjLmRs2siykd4s9BMXLIUqN00BH1sZgCYaM/i
J7qYXzVpePYC0dJk22CiD2sjKjNsDjKvyuCoMXmfeFl+ByyG0XJUZOXPAFnxJkHKI9c9e6DEziNH
Ml46dhFC2PrXzx6BA3D8T6c0ruOP7wWQT8mxUXHYGpUxYwiZiZlIB8WG2OPwfGjf5dIxT5Dl6VqW
IaBC1gshArSNh0S5K01diqfJglYsD7sDTf8zjrV3qkUjUi3xP3poylfyBGCSlEWltNHcVrke0WWu
wt5+P4vbCREswGygm28tmthVhqI+a0ijcMBI39dPHjXuFzXl6uypTsaCh7s8GUAFC9S08mV0bBdL
hGxd0+Q3RREu1McmyoFDhAhDf588hsSlR3y8JUw9ZlwiUl/cq5U67hRgyHe/kAhAlfVXeHz9z/A8
ZPYZUcRt+8emAirMQif4Tsas4R4Pc1pS9BV7ZbMSp6GAsB/UjnLSl4BZaAFe+XuolS8BEOkndosz
fttBthck2pK2VlCnrvnTKx129GWYzXX7O9aKtjQ/ofoOnXVSIwe8Bqur0KpjCO+SBwHBct8dWyp0
fY4EkxAAGPeFn153zEluEdNff29ToBIEJ7Fh3QuYFro9QAEzhA7giNWkKrGO/zWWOx4k1mO2a55k
bJwECpCO6qTWtxABig62GRyY6p/IQLcEFXDbD9NdzTIDKmRExuajPhpKqTj0jg/Nad3bGiwVv1e0
7mnbkiaUXpCXwR+3Uy783X/y3CyzGjGYzUllU/lFTC/ZO66fHKb3RL/x2FcnIIXuzhY3MAvjlNbc
hq+1ZVFzR/GU7Gxp1B3whEHb19U9h4w1NZ6T9qZ9RcL/jKMmJlo1hQFiosn4GjruPu4tiDThxMh5
OUAUPBuq/+1MZ0dH2HvCkSI0scm915tMmUSVEJ7RoR1HiY/jd8T0kM5tgPou3CTv19VqGwOKU3S0
q/XkiY7VITW5qgNPOEddvsKlioIy/QvIjgVdV3RW4rKdqWXx0ZkegkwCwXE6OCG9GOPNtes3CUEV
cHzkYAAaaFh6qWRwWZUR9b2oHmH5Ps0TSkzZrQWWOJ0j4M2EgrYpmWieybuRWIWk1W2Wmuuq9DIp
wQsUgJdNOvL1rmjom9hsnL3FKX7zdDn4S9ozuQdYtvfEHr0AcrCBoMkXB0wHTVFgEPxNgiYijV97
qrxbHZH8tgDAF2qstOy9rC5yjwLXmomuqYu6GH6ck371fa4eOf8N0x7lUMwUTjkOGe9MZ8zD2pk4
+GSwCthIEqlTNDiq9ejkEh5NFBKiM32kJBselzHm4cI55zP9zmFhF/lRFiUnHVW6JaczCmxOI8LK
flGby8Wv6yMyGRC4+ymCtRINAFfygvKqJg902sYsgEl/Tbo7cIrJBo3MNHCIylM+2sW3fRXuQ9CH
nVdBC07xx1EPEphse4BWMuK9jHDp9rjcbgNCwUaf4uJmMBddNNcxwOkNwR/ySTlSiN23k15IxeoB
l6Z1MY834PyQzu0xWv3ZekrrIFBFdvdAW7NhsSo9CCKYuDKayCCW04uy3NlJiUwdT93+eQKEJbDG
J9Y9jEehKJGshSK6evs4pIH8a1YC0Jc9uhG/oJuzIHLdJpA9LMl4Rl3rY4fLG+Rg5TGFcOVllARK
BIvfpd+/zR+QhhgM5dufu8hrJKjRybEQKDA7MNRYMfYVeWuKidLnvZdggx+wwmq4AtddYXos+hkV
9qor9JApdMPDbMb/ifdfkzqRbo17jWK14nnFvGBjGLoafCHY/NEeR0zDquNtRe8D496YV8E4+OnX
xb+HCoSP9R+BqkfdFtWxHZuV+poKNlpsiDtXjF6IHw7RpVEOFOyXb24Dcb4P8+8ln7CsFibrRApG
eZRDtILLuU9d35uYxfEOW4u6S7oZA3f5wgsM4MLepnMz8YeBAJzpcTHeDRcxmYBvz2sSmqrQaRd0
IJlS8Hx6v2pwrVM5wBD5NEQHqaaT19tgzD9DytoAZUCjzXmMoSfB0KKiscdO7mbKrA344JLwfXi8
O/XgmocDNc7Egr7ztjPw7PAUsgn2+q4LW4zhn9jTllAlsfKKxUdZkdi/KvBd+s9R3EGF5POIbKq8
cOsO4AJN6o2/KQ1WFu+tcQmWJUKOHajCVOoIsxLOr7Piek38F9nzjkr35R4HtxBS50QDW9ZPXPmW
3XRTb+wNU8Jzz9Zm0BpqP4h85yr8qEoEGScoyjtbYPIfMedgNTFkhfArTZ7yPLNxukxSAwfTPYjC
5AO1i/13gGCOE4OwAqc3+fkX63m+HrAs8gP28e/VwQA75QrAgFFIMHCqWpepji2duRpKB9RC0YV8
FeqNIau6pygpJKPX37V52HosNDxbT7TYDEOwjmRQVjMkthwNj6FuymShdx80sV/QV/Q9quXiHTTo
flp5PDkqslUunDJ+whQoEwwX1BtKcWpLzLJM7sCkOiG42Rd8XX2zjS768pYeaWH6B02weokbJfOa
a0eEWWUXUcbUgzAzHiptiL+mYrzM4virGxi/82tz8bEaxLHr8f5pOBB6Y6RVxAie+OEWr7JSAiqO
GVTfUbgYpKmdUDHEXQbkhUNz3tfCv1LvFvRf2SEfLpEpyJQgJbod6lnb74jCoDlFjkmMIccKLZ0m
+PQUvVEF+aHpReBDJQsjMYhl8NknKE82ryZQLjqCNat8OY0sqSZfH4vxSi0jlEkN4O/4t+bxYHFp
duRNPFvq4qjbD4n2jxarr1C4QhT/3pPdYSqwZ6i0E6BedBzv/QVeHe34MvZNCbbEIvMIl6VX8L3M
J/Hnf86Yx+f+0mMrw9tKuoPcrvdhCS/iOBz4F5fS9YU38mWPwKa80UixxE6k2qgOktMz9GqbKvhi
nEBvlIjkQBZJjWvyDrgmcvxaaVOTp2kUCY5Taf7nIDwRdSeG/fj7QZPASgbDdBK359B8LqKsmYWB
6CxuvUcm2BVqYJvlz6O/Ty7//ZrfCNkgSpXP1yH+nz73itc4WDfCcw32sfhPVHs0w8XWc9NYXOPg
WBZ982Mp/CvaNkLP6i197/0f8+Oi0+yGz2jfFPttAWvSG7elevCRFV8igJ5c9M9FIvwaF/+AnUXg
7PgGrOkWM/4qWitafehya6lHVU6GEb6mnE2nyYNglObQakS0nnw4kOXFJB/hBEU0XZz/SeAp9ihZ
GfopcZ7QQM7pmul8lwuwdMBRcQXifisV4cGxbcogyyWF7iIJ2kEEQ5ypHGazN9T3WRc1aA+Y5gUG
3T6FBsZja+hXzXM0UhTHmV9x7LIYCtcReL7kwl2jyUSs5+3AKL506yMX92YCw1EQXnUVcrN8QALF
hnheYWrD0qL+gMOowBKkIruX7dCJLb+D1/WsymU+LxoDcldUDxV45NERBQ3hjYgV8lLljIIVBXKX
zQ3lKMTuEzEdOmQ+WaLEMU4VI0VALmSUXoCpi03Tvea9btxe/h3Am04rtBHlfzo8mJ6ht8LEgzWi
GlnbZdApFf5svCJaE5Y5ZLub7k49rBtEJ58VLfCCEsR4ha6XsZSS5iyVbbxQqr2LMruHkgjAFYYy
KthkZ+d6Hh6gU8JkGk20P8DTsIi4i7z63eCUHi2lugc/XCw3wRenRGwF1oxTzuzIdpOv6R9o3RE3
Nx0ehOk4AjS5m7dftUALJZoQj2EGoXpnMWAxyUEY87zZa5YDaOjaujiW9O5uuL+gLtCmazLXSVtI
52l+peS1WCQzkUcwD8tr0Ow08Xzh8Bz4fBMvY2YAIMzZbXV2A0Cirqom23sF3t+OZfSrXKD9+5Gh
sJLpe0k1chNqxJGJP6bAMQghkBgDfMBO241La2bYIe/mdrY+W/lh2PVag464iesm+mCZNXLWbmRr
oFskqGvgxM8I69zrX9m+IP0NvO/IIbI9NBqHvD1JLjiS0uDJlP/pHX5qcoFh636ChVIvwpvzcdYo
bHboyvStXZS7TMOwWq0pQemvKEY7TTTNxYkLvqu6GKO3rWJ+KQJAMkZ/vI+6Z44sM/V4/46VWgVv
nAZOu9Im9wiZgbr0hFGoZnAV4eZVOG67lVum8ZjBaO//EXRKUvPlwTwwdoxJ8pya1F7/WwgDKi16
QkDTRly69RAQyNnhDX+JUwbffqceYcmzLmf9gO0eHFhg2hsuVvPfff2LYmvdSfpNsPs5XOa5G9GY
BQjBd130hMK3qsmCX7W/xBeeQbl5Or1gNupXAkm6xI/BCJvb8Vf6EzgmTs2BlcrwasBeJF0h57kY
0fMJa5qu4xSiiveTbGNFEUP5w7PXssswy5eHwK3V2Dj0LKq2cPlDkWK573F83wTTgYQgoBcUhYWP
y7SO/e4LLxg25QRJiQOVdWwH2w/dJJ1e2jMK1aKAzArQEncn+mZOBNGJTbkrl1uf5dV44GtrKc1t
orjuZhZwdT79n27Zk52mkNQWLBy5HnckTpuMwdW3U895l3d/km5qwR1zJzsTdRBj5yOWIvkjbt8R
+x+wFwFRW5z9OHcZwK+sCozE4sLUgPtsxJCY8bdKh9lkMI0Tu2BXtwxGeNhF6KcAB2o8ZlTAgKi0
Mp7vThZJxedEio/0eEd/8ekWSFj+4pCpwm4r6YqXirHKlHPbqiUFdvt1K+J1/vz3rk9Ouqw6Y9+U
EQesxhF2coEqk17y2dCU5810sM8F+3bIdxzN77M/sLQ/954h943UGY8j4Uva+dePSBvIpTK32wCz
LtjSMbZiADzOGUMKanMmdJXSst04vN0sAVIeWpRypO4RlDWmUaZaAMPjbLe9trXXJc/N/l9za2Ma
tWFF9CSP+VYP3EzKmCzD6zFPJXD4ec+pwqAYb4xG4x4XV3g48F9O6lb3pm43oSdjmEcC4rc+ppi9
sHFrU77y3lLwTMTjOmpFuRSf4rBaBoHawo2XEpWd2UVHiT45ri1w6zwKHmAsik+e8fAX/kSibdYx
9l9dHgjd9FMXL5Pw7qFWA+LbZcfT4eiCSBUt1f6Ue7+v1KqN6qp3v4PNh/C4zmpxZtkhYiuotoKN
Ub8p+C0vjwD8np43/N0AgzvOKby42+Q/4xNfsMk1eoTaGfLM4UpN7Uz6MDqB8XUFRCndsKYkKWqf
7qkjjB/FrfExxGN8zouRv7tN1DKjg0iUq5ng5lKxp6XubUEWsrydqEDgVXz8uqQ1JjV6+6Ah2Tjk
DWUyWxMRXsXArqKlIf53mTuHW2UtxO75wxShWzFVBS8tFuZVogLXy6+bBGkZ9QjSppmxxHI9jhTt
MrHc3HW72zI1+Rb9XAGyF8M/fE0x98P3UYzUD6QLik46xejZibIU1zqx5hPan/soiOguyO3lCuA8
0luAaadAQv5qk6Dnk/5hXcjhlLp3hhmets7DLeAk8ghif0HmMpjO+nxgpaR7V4+2FFoGPHLoaybL
KwHPvzY5WgUDASWOVDvXdMJzmSuu1GwtkyzpHN5Pbq4nxc5ZM1y6WF2zq/dQFSlTQ4DOjWG7Pm+Q
NzsrFd3yQsoVWOw6Q+WZ5ishVbIDBm9NUo1MS79sggPa2M3o6MbkiBPzVQjjvmpDyKwdXqq7t1eH
cJ7cDimuyJS1abKDM3miwgss/aBm039Ik9tM9X5lIwLEtknJ9N2gS31oLbhTKBKerKGL0jcK38Mr
I5okKIFjiZ+IzA609M8UpEfinJ2xkEkdhpJ/160btooVaoMQtBG0T16Rs9xHYerWV4dX+0rOl8Cw
ktP5ITh0n0ywOsyMhfIcQfu64AlIwVYBXkDwwci3NeUuBf12sAomERfzXJaNJeJYeAnWgRJtB8cS
bXWS0FH+b3rpTkrBvuoY2TkhQQ4fIV5OpPe4Q3l4NPzfZ9lqdmuz1nWM33Q9QCWMv2EVRrtAIt5U
c/3qOgSrdu74w1epqeSR56fiKhv+iApAtQPa/HWju7l3PhcHBQttjnBwXZqdKXO7MfpNvZhISGUQ
I/GwzHNNs2Kf0IQ+aVLmmFrEZ+gctQrkRX0Qmq+cV+F2yzYr9m96CDSUixTp2+krleyzEaA/zzcd
JPnCS7DZn6hWM+iGeckZk7GmnWBnDABfnPjs389pCqUcygO2AG60Fu6RCVg6+yQeYk5d9arlAm4d
fZXATmYonbjgPLDA+BzJiJLFgp6hgVJEO1sOKcTvrhTD3xY+6lcG+jKRgnJKBYxAvq0ytuap4bsQ
PZxG1Gge4/MYH+KnZVYrN2utnL3Z8Sb4i6DEfYyhJm/0SnxPom6IMUhovHDtdeNoI22tQb4vx1Pf
AfpKlO2m5lSEYozfi4aHga7cpGQxtRh3hPhFgWD4q/lyEOk2DsHfrbAsFzz6LQjY563rRL6DZOrk
VU4FJY+rE8Lu1U2C3UDDr4eBscYHMmCxCPXu2NXjz03DklIz7xm8Wt+U3zyIr2Xrwqjb5pAmgrPP
TdaSejZeXtTBKysIwtdDjp5B6Oq2/ylHn6OSf5tk93p8MG2LRFCrabzt4Caggqh5Hb7rQCV9v+Ou
Ua62DV1HMxsxFsy0kArHtssKVhOLucrIkzAquhmTZkTJKoXxqdledNicxBmQ7ONs0KgKmoDpcrjV
ViFN5WrcLzRh7Z6LXdnykOUfcUCuABOzdv+9DdJgSEsmHvILYf8RJrpJnWxy90AqlrkXMsGIf8rq
pEPDI90+Z2uKr6W+0tU2JPdoJVpcXrToHZdxMzBglr9RrLDIcaIOQAcN8ohEHsiPsEYb0pV8UEbC
SFVICiyjiG5V2EPIVKQ8VfXsKR3LmVUTF8+hTiv5PSVVACkeZq63C5v/qQrP71QJL0VazTMb2HD/
tqMNplMZOulyJgUjLMWgtQhNXXTE9OBOcKjc1xAJVfWWEQ1wlNLCE8+Z5Vdo6T8TsgakNmLdxrbi
RfzAs1nuURIASKcx2BHmnLiEdoA/Ifpx+LQLOBlhWHLzkLD2jlqoz5ZIPCSk8/i3ezcaNyrrm58S
Zt3qiXcfC2m+6JRr+JXRIpA3KYgSc7zRj7N46L5sOb7tzoxISAu6NwjSN04hG/iW4dA4yE5ms+0/
OBOBdUOdd6GJj0XZk0EB2eqcSg4uI4rb7udQ/wk9nIBx9zjEYJFmZ6Fd2YsUH8QQ6CWXN79uWjyy
3YIhKL/c9eVNaVtaUwyXCiDzgMV8dCQE15Mj4YpfT5PVsK26yEJ6h/7NFUD2VHwy3NKtulKYvBzB
uMySDTKwKtY8aj6Em8vYSBNfPSvs3Kbi31p/1iWMJQuYEtGjy4C12CcvbiV9rVV+AQQVPV6n5q7j
dCsuraOMWeMd8lOiVqqtApJ8C4ZWZ7q5zrXF2zHBmWQm7uPTFr4ZkEAWLQqbv56GU5hdfiGC/eef
gtMh/3BZxaW4EZMRtFdIt8klzimB8H+7eLRWboUzcGqc9KlKRki+F+mIPFlYK5ELcZyPdxP5Jush
jy+OM90Y+CP8Iijuo2tUaJ8iBuGz1lA/QkUiXiFjji8fSlDfAC3z8wzI38HEOeIePxlCkYEfbnMk
s2V/siakUEPsDoZ0VdTJ15idnJDNnb38TQHBxs8bNKpxaxFRq3S1G2Ytd5WEtfX0UnikA15EWzEf
apcXAsEQ1BX9U8UtS4hv9SSAdCbX8rUPf3lWd3tr1FAwhSHL7fHhf/0YHnHLoS3sMeSz0gtdRSo+
HjpRGLkvdsUt4E//jWWqjG9fvJILrnE9hhSiMFl0CfLsvSzdsLuv/wQ0Xe0bfwtGxGn3di7Q9Kk7
khzC/sEbThETX7MIP8utfoUEHmIzLvahwYoXDZbwx+J8OIbz1GSKA85AOqiy00WVrwa05yirA4hp
y41Kwp7VsEvDKKoesJ4fShRAuzpc+mEMV2Gk4EXbKL39EvBQ5j5UNa5fZEuAceHZNQVIayFboRv4
x5ez6M3brtXkcylOe9qJsOVhLxC4tp+eDH4xQi/Axg3xpYI4QgX/IW0nRz/g3+YXoPNLy8oXJAOt
2KTZZzcF5tGckmy8CdNhXG3BShw50+ecpUr8XrL9Lpv+ROCixEhOiXT8VdTl5CGHx4sRA8dYtMrM
wnC3YJQvxcexFqq1a2BbIejuQGSOXKgtN0WUUiffKyuvRZnhgIVoBR3MHKm71TBLNTgks7J3fjg+
rmXBubqJq2ZEKILSqq5420dnzl6/wz5ZeaxmDvRZP2TXgnpCZjWPAknLk9CMC2t8PzNsRMJdWmB6
D91tABpqVySyEiSUpzQ9kamxnpLCV8p/JBQCwRmMtw+9wFRsSYIsKbbfkw/Ik4wrem4gWkcGS2X2
IYyDzJLnZrbFAyUs9qttZJbeNUhLolrpwl/4h8h64QWIE2uH/FSyIH+oj44ADsyjyuPINWILFuBC
HMJxHxsWX5gRurTcY144UTWRkSMqZMuQGhmTKQcK/v0oDzXgfBMoMmVjumTa0jgOGMR9C8IzXuVy
aov7dQyxm6s/qkZ93aqYmxdAOgHVZ2d++YfeiWjdiW7xEbGrFrK2CHiIMcPgSJQ20ZaWCDlar9Sa
YpIsbb0e/Q9shFknM6DlycK6G2T5Xjy4HbXjvdpOVzle9NuYSY8vC9dOcc9Qu7gH1HbAKLGeuWz4
ODTbGLevxPXKOTTJCfeAo5r5HEFUo3GAUzYRKGeiJK6SW9GFruayR97pM6Y+Xq6/+g3h0XwU55UC
k8HgnmL4IsiDeYihRwGZEYoc3Cb3Yvc6sMKmhKhJUXRKTyOKA83m5nTzupUxs54J+kED5EOzDTQy
RQsOoROxGKVjVFbClPEaPUNqgiIJEl1lq7KDhxwyDTO6BRBwQx5u8Xd+qgGIL6Bbh/VoCscWr8kj
jLSNRl5FAtRXhQIM8X4E4hyjvtDY0ddGCKQwp9limg3JT0v6Zb0Pi/nmeLH4cEoh9W08rssxTv8L
xkUdJ0cjLnVIxt5RrHnWuVsBIQ2QGjfmEEwl0rN7YFW/HxTThRSwJI1e58TSBoLhlrDDsEanu7Ua
fkD+72VQUxc4qZZaFgOYUJHOD76sZ3SXL7Hw7D9WlBYryMcPnAv74hvkw4D0Etu2Yy5MxOhJo5VK
Rsi2i6OaXYgb0ev+4aLKEbzbdUHANvdoEPE1lwj4iUc7jL0fiz25thO/r7nuBHOe4bk7PSzFX63W
Yx1RD0iGBefEEig0XbxxNRdh4hgb4t2Cy3ThvkkMZscsvhTaOd6G/nHnh/qCva51c3aeBS6x4o3p
qwjEml5rRtw39HT1/ul7nt83S2XKgI2X8zAftf+RTYyCMH4nlCkcqlP7jfdzEas5gnJnKA8B1T6C
ZCHvnn+Ef1pU6fCxD5DFFfm1hDz9tDZmRKeXdE0/YS1Zi4+qH0Zrszm6c0n2B2MWGA/o1HdfklDR
YQSrtJMKQ6iZIsY4/wCauKF1XC9A0+oBpq8Z7fHAM05DfmYcOVBNNya6GXSHHha835Z/NmsHL7GW
FnAcoFlNjBj9Oi9sGd5DdZ9VVcp9wcFBpojFcz2WKjJ15dVoEd3f2Mig7MBhxeaMY8c6f9OGHQ9A
OjdqR8XHs3BAwlKPNdmwSSl8+lUj1SIUZPIGJS+c5I2aavZ8DS4+bLXlCvlphX1J8zNhWMFtZWzq
U/xNo0Z7U4llDOE+sm5eO/tyE1jhGdF9Gq5MoiC8RCDLttqwwrWU7UvFvqfc7c9KOIMJW9CsCpWt
kTlU1YydQI+9v4JzaKaVB3ClSEjzp+aNzTNcUQzUK5BzAEW19IEEBbaku7KDhJDlRh1Jn5MzlQhC
bmgbYW6E6cGqlLNqBOVdhVWx2C81DUAyRp+4mQsv1obksUEuMBwh47rqkKkhEx/rnA2P2MQa047t
VDA2cMApl/7T1e2dVog7nChx4eSyZO4GWZvNP7ooL2GBM3cwAArr+hd93ZUPORlPVwMHiA0NuvZs
R+i+Jt0l036BStT2G2xDCL6e1fzDT7W83pcw+cZavhG+PoNJCDKEtE3wMoa03L5Vy0CN1bbgDamI
ADXfMeQ1PVj9+dDvL6Jd/0LuJnkcgjislZ1tYrOmH11DNDz65Zilb/XS6P5CyaKhPahN+1XGJBZH
yp4HO6H+ep1RO7vP63ibDZQTSBUcokWHSWNJA3lLUZefMVgVpEomi65YZmMpzLZ9+PMkskGwCLFw
j0hJpAXlIit7PAXyIk73GXpXf+0Oy9X3cJMpWj5xa2zwboi/IMwQgzTYI3ISkQrZfXCQ0wz+dM1N
hhPtATk7TaRfevDQup3/HjttMqaJoPRdEYAXUqA+gMK5r7yfMISy7oBkKx8F0u+LPXcUJgVjhX/p
YrotuizPAWg/Ofp2U4O9r3X5zw28oIXYuYmCWf3+4N8pvMErYSStGuexMc5+rvgU9exLZvYmkT0D
qNiXBCsQSklox6ZZc9UgLUmfgT23Z1TafDv4qSF1K+e5Vrlae52nQbJ3F5baCRWXBrY7KSJ8H5iz
kkRmeFXpd+WnXcmdun8VwheNaN8oT1syPNz/vMnKs9HD7g8XKiL2f/wgbSCf8oxfvQ7qUtoUQHMa
E+K45kcWceTHgqn52+oIwdrBlxkbXAQMBVSwmIvjs0PBQgs5MAWGD05UkFPccpu64nvWZrHcwJHN
AjYsN54r+QlGjZvXRIaYQ6AL9iGS9L1xnGqIirp2Ou06P+crLx1585lXHqjxXMqfK5+WMsTdpxI5
BlJOfjQpTUvLEvfTbKn52r0U5sTG633F1ehy/1lCKJJpbycE9TIveG3aa40i3twLUXiwDxSu/ZC+
o+BURnATHYrt95KPsQbJ/9+1AtIsSwzHiSnWfcVLV/flLGA8iCaND+gTaeAt/WhfcEAeyqPoTC4a
tFrClMmu3KwT7u7mhUMK38LPFtyHNspNAcRy8vUZIZ7LwIjJgfIHpxyPo55U+59bH9lKFo7YbQAj
3yCaxABuRBmU1J8PUySXLTxNpkCQaUooe5n5AHMny0JnrGpjbZnLcrk5Ep4ey1Sp3sBnndYP9xZK
s1d8xdaAyUxTnok7ol0ZAOg7QXvkdpuVOdXppy1xvrvEFUrKhR6vKBIDI6T0dAoHaAquEgAIncYb
mkcbNacJ6uy821j2C2na91yFk6NiMs7FOf3dlwfkFxtbERP+MXX7sIIz4HwdJJtU1TlKkPTSO590
h73gCHlyatttpfVe3Y2fmQ5+doFeDg1g5q4dROnPPEbLSnbDPhZW+l43EObg6YdcggRn2BzGTIMA
TErw6wvJ8aVPL41Oy/CSY8APhXvCcxfEjWdmGJ+Tyoe+Gswh1codEJaxsDwrsPVWcZx7jnckzhyB
BYboUfgfif4GaJTSo1tQmYh680wlPY2/7/7gJ2BhwiseKfDyNexYO50jhHTuToSqwHreXNVjUw2n
aJlf9bpK3eOUXrVjvdBk+9X7j27Wpa3QJqlLxDccEGP8wUER/iR5aal3Pz9EaXEg6gf13G2dkmaP
VoEDjO1qIhlzZIgOBnYxlT5YeD4+Vt12s1fcXzFSZP+ZBp5EZ/2oeCEQxmeodCR1vUAlCmFffzHT
q8YkiBaDaxcGHuNte9AfS6eXrYWOb58q/7BYFGaPqY/QEw1IYCuJ4dQuWROUuHDikgC1VTvtF6/c
b1DfE25OW0vQybzhIgpOFxK/7fbsezs2XLUUtovhm5MkNJZuJGDxh1aOgmxpmp93JpAtKyWmZn6G
i8AhH8Yg5SW/17jZp8jmDuZYtBuVq8KctBeqsZK7iws9pgmwBoFj1h3XOtGL8D92GSH0PUCLKLst
UDWPdv8Mrs9p+bNa4Ms8zvH2Kc+KPUyWJGkVF/MSAGf6xjf68AQbPOktyoUeIC/R91mdKEIhck0o
gcivr1ZE2xPufETNZIctSxUlHhEcG3drfRmAG9NAmY9mTa8renJDj6Z60eDS+oiTNT7GEPHEgdqI
YbABll0L8W2K1TNbPdaTGvQyX7KJ/vjOsZ9lySDfAFFJiJjZyql94Y/zVdMjZzosWwPvBen7A6F5
zigC7gmyYRsmZwWLFxcEi642dfsseMXyRbYqgDlcNiDmqD4nS2SWbYvDq/SPLRacaLbmgZTxYrla
cOfh8cJQMTFgd5nTQW2WaX3e1/L1lSMPIthawAE0HxOWCxALihzyS9DiYw2Azhd634Mxj4SwWKwn
q2FWfamj/Hn7BAqlR1anxhfEeZlsmbNhF/ePt5UHtXOlQtIEtQbQPrQpUc0o8UI0xnIvN/HT4tVJ
B53ug51VYm9aoumnv7pOCdhcJGexLzaxVwm+X25Xwdq4e7KVd+xGnRRjjq5ATkqEcMgQ7GTUhMO2
pz2HYpXANQJTKwloX525rzG0RxByjEyK3X7paQUxiWt31swZlItgPPq/TYlREGcpXoyWssARMDxq
G4lmG5uUb8IsRfQbhpd/2fKVTGvP8DQyH4pqJHRl+ieKtwjsLH46NMQ9KAeeD5PO110MH7C6ULBl
fN2Pym0eVCowFGTETSTEiwDnHWke873NMXHqrfe+GANGu7dlLfZQ9UU4K7NdK+bnDWsUVlUJAimB
a0ltZXgpBo3aN+w3GUJnpBASXQ+dGDWa5lFo1DQa6NDESrkQq2CiPsLRTdzoy+sUP/hni7RGkKyV
eODY3fz5jvdDlGLWLwMu02KB0vDl5x2k+FIc/lBrEN34K1PkP2B3CqJdiFnS1p3NJZBEjtV+EOcE
zTTpp93jacLA+P9sFtfJ1hgCdSfKH5g6w+1AL2PIc11k/gWJBQmftovZqG5ppA3VlIl1xrlGRbNw
g0M9FmbM4oNU/mHLABtqD4iVzXA+zIeeSZyPslbLfmvhhCjA2m4lFjxvpI5ziyvpKWwC8BQehqRu
70ilG6ii5bFIzdG9H84vXQqHoPvgxeWF7nNlOQMumP1pR3rSfT2qgJw04b8+R9jst++Z/Gq+vjeD
gL/SRa7Oxe3fzK7tqOIsU55g7spj7Ed2gmv5Hkv4GQxEpuP8Kv0es+FL+OwUA9UWTLrEjt3uFyrV
jvv8QyllTcNRogklQ95O0zjXVAlKdxLzGFYaMBMzyv1CE3wqDo3e+NznV7zAvix4VVzpcjDaPHzq
wIe5aksQoVqzEN6RwHfqgO3D0xrwFtHcKTv4NKUpMjM5AdHyDUUKIfhJmN6Pn1bIruqR9v2ZXFr9
SRtc9kqh7JDb9RVUMc22EaTJ27Kxel6Jla/xbjKOPi9E55vcd6JXPAialvP7UFdv+zuXRNXRiFwq
7EibGDNCXqx22MG0uFQWI9lufjS3nW/PeaVpykt0tr6YUXfKE9ZzlrmHRzFRQSVqb5quls+14KZS
gJzVoTRpvhL9zxoguaYf4r3QxMmfa89xaqIXdkVVDOKxA66nwN+sFXS9abN/7Aooar67E50A8GZQ
o5rSg7izpZ4+xrn8xrViA3HYK73fzdlecw3ALrLhR5x5SJlEXgSj6mvLWUaLhNDpALYo9lB2jfz/
939aNn2qzsJ9WyDFX2GYDgi++lTgpirfeGJKA+A+CJK5SHdsVslUzeA+oCAA0i371QY8lrgodL7w
yKxlUv0V88BvHADVPem6wl3X+oHSRVyD15RCsRwdQzAe3aKnz4INKBhlhGi1Gz5WuCHfIRamDASl
OLPe3XSIiKglYVOx5oeqyyGHsu3Tfj3zuBjDcwWSFQO6oxFSxPGdz8IHKaRZlfuniXt+D3cbKkQ2
WF4UUSEhurvlqzmGHuhJ2uoqk1+RQMnbBFvUipyUNwv5qYqzFUvllKnxh4Px5ZUgPIt9nwssgKLd
hEJ9rI2RplQzlAu9SthA6o6Y+9VsCg3dHsVoc7UHjsJROdAqVY1kHyIrTgr4Ng9NWQvtGiCoXZug
cmH8HwI13Cxvu2x+DxTTzq4CVcCtVdqPr9+2HYY6dYZ392q+HDp5Vu79j59RvDX+tWfkHGNk+/M6
N5TYLWfmDt+wpA4SxZpjm9Amv5pAJHuKKxZXKvETH8b20LAv1dMMilQ1l4MTBtTSn7O8KKAz+n/c
yZTXyugT1PGmCTWODXCmjEdWsPgrgE1Pm4N+BingRfcKi2jr1IsSSTxCKBKSNzT3Eql8C2lPlNMA
CewGa9siJmSMXKnIluB+tjUppPbjlWQ/79U/4ydGcnyKHdLp+WEwJD+zXIxzE5B+Q3GB7K6Gp5rt
fpnJvZZpf3AANox7WD9dwVEXXSwAYbpnQektGjIdUKR+0gqu1uo0qScHRMRR2HZx0iAsV/3lV9wz
oMmx073ktq4HCfXI2Q+oNeyx9ctW/cabmBUqNVFmDeS7DqUjQWPxICANdXW+UWA8Ht29eKW9RH5X
flJgiDVT/pCWM6z4t8UwbnUy5ax1yOOSEqNnQ//v7IcCrSz1Tr4X6p42QebGskEMKeK9xQHg5O+E
D3U2q2y+aFUt3bka2Y9XY6lp5EvHML9Ro2qqBgAeKHXpIZO/IEkrlH1S5UDp1Eozt5Lh2wnZHJVM
nG0WzZqE+yteN7RGHoLZvxHARO4VnGcthBxEa5idDKB5QvzdKsa56vjWS0WpLN8bt/g4hdhRL20l
9UJsi5M6ZbNqgh7LnIzz0zpUAshx7l9HOzhNhSkv5mymZ6I9aK9SQa1LBEEu73fuFlCdB6MUhnVJ
huaTl6IQg7eVVA/n1E6TK6u4q9OIiblM91I9PSomROzTyU3x/W/VOffBgjZ6jOsdXrDS3zl29uSf
Jkqqw+LeAkazY5ZUlSoYNoCWZP68wFPXEKajgI48lCyDKAMFBpEf2UEwbNXEtQ8LJiB29pddnigN
6jyig4E664REWmwtujBfEB7XG71d5YHbr6NqsaZQtjDP02M/Bj5/zaDx4WvwPv1FM/YoYITlAxxe
iBkIMXsfP+IY6fFRo0LOq9LjWMArTvJDAy/0ucHcL/oTlkVagZ3GmvqquOlQ71gGFfKBP3VnGGN8
dRhFnyEqtDIZrkJveAm2kpZHPz4W4LEY5rgP8XynvKNolLiW8UFpycCIZAILn9HxEpHWDW/aZSif
kMkIegqnxeqZNGHOL6+Wf+N+fbO1ALXvRklZ+FMkTmG5XoUBhpWwzaBoH0/pX75x23tQ2XzcuYUb
tVR5B7k4jJy0LgbgaFCycjg0e/zSbexOa3LIzCqyV9Lvf5WfvlZnVFgzNUW6R8a84BEb7AxIyF/o
v2iQrz4MXkVzlV+gfkSDb2JMqwWT4iMSyBTQ6TyN0TEwGNu+pCN8frThQYa6S1I3Bf7u15C5JKjG
6HglotFCGbe08eaNIazDT+Rh9XEWBFuStMlqtCiwq1GLOSCqN38plOo2+rLD8kBi8Aba08b2XBfH
FRqlP8BM+2thfh4oa+8e0WPd5A+TnDM0STLtxOmWnKZvw/S5sMc5kGzt2IIoNiZzNJ7mly3CgDUy
nN82OfF/KasLtL/3h3G9Xj6ikKc1NVeTy9pzq7P/YVTDwmdb930ozyVbGVu9dSCe2RoH7PCf+h7Y
OwGGMUNwdhfsNx+jBNUIZl2LNkt0NthoDgiknPzpTBWUnstDwTd7Lapc7jia3ZqAdyYHUefKHUOr
488SzCHg0QvOsOXnWuwqZq9SDv9v0z24Qjk4hw6qOzvYZBf9W5Uf4oLk65ks8In/OZlEUb64vsGh
XdhXl/r0owKUB02lJyCaDph+Mb37xqZWAAwZVMJEUo6sQTVu7G/nDxO1pMkG+k/9sWCvn4JXVE5B
cYlTPZjnx03UqhgCfyGfsjCgGdBfFOHuWqes7EN6lfsVCOnRPOBqa5payyJeJbwxKddjaOV1ATft
Tue47IltvRpZ+T+zlZLSnUu8coycCGyRbWu79xoEX/WWwez+NzW4asZa8w4W0J2MISUTf9mD1Atn
BZ1IWednfiHYjuIvxzyckt+s9T2UyHkcVVRFc5dv/q64B3VAqWKJa8XiuZS4W/ZM7aM5jJ8hhn+h
9Tg2YtUAtSpaz79w2gu8KhWopbqjPgWUGCLbAKOCsi58hL5UeOlAXAnL+Dnh7zq+BcoM1WfdX/bR
d0zMb1+Rk8sZE8tzQwxQhIszIIyUtmm2mpNls8zzBSiixKj8Zpf30kISHqKZsDVeoN4DegGNj/D3
JTW0Eykkbxrnq662xf+LLxYD4BW8f5Ip2CYu0KaJGqUl1WuIkzwxBC9lfXGiMNduggTmmX03yHRw
ZbLirKA18g7/us5igY6nKlEOaTb4haHEXMHEBvliNyq8le7dkqDmnIzBKu9b2kOKq84G9LjVeu/s
VrExDwanjBrj4o95Jplr5NL6F9xYmyznkfwsrVHwPSOo93rsyqpCY3jxiI88pMsrpxq6bAcwxMFo
hcHMzgcHQdbXV/3KbszXO0G9jX0p8LUadmo9Jtc/D3Dw4fW3qbvzedY67Mtl8nRCVW6ELZ/ILqbM
7obFvfFhv9+a0Pgn+a3Ue7bAoKzXJ0Nu/4vu7cqb+1eWub41Kb7Y6rISiWqMPfXv7nvZIh5FzK7x
6X/umeX2d1pAz3RQNXhL0HL+slLEJS1SD6jXF1VOBht5vz7zCFRRcneqQy5EzPmyfHmD3fhMV6ob
s5ByLzQeebAof44UjzbTp0wCBzThFvqkn0blSUdEx3Te6X0WMtzfEpJ86qOh51gwsWrGsf52+wnv
iZbOpekTBNoWJTsJYGgORgsXj3YoW6R4ZGihMEJmCVpDsFQqjjBnMsLROUgLuQJrg7clJ75meC2Q
oMofnH7qyZ8p6WjNFo9R5tDm1Ip+/TbeRNWkbnP6M/CthwPp5Y0latksIvpaPmMN5+mecJA7nlp9
dSpjeKxBvdArukao+oHq5azn3mcC/LLZE5EEBSvnss9XawbkeHDbk28pncyjzAjnhSAPQPB2QpO3
6WkY0Upz0WKl5im9r5rJ6Fsyz/naT2hbyW3/k/YtxoKrI/ZUMEdr4Uo3iMWC8xTe01HQUxkIrUE0
mQCc2a2uP9uiU0Y9Q9raqcUkZva8dhD1kV7Urk1DHLWLbYaq64+WuEwMIxKdzKPDCAuBR/CdWxN3
awhrVWz8tHOXuUC+utvFBjtSB0BWKOnjsKK2HpqQTM1sQU5WmI3/bmL7q8QqOjnhZRDrWRArfp7L
HYbi7Ys3xykgFiGBBbvss4d+oL9jLPhrtpkeQosqfha4VNFnO70LsOwEjqTf3JKUAWOEXqGv7Ff7
Lt3wHTwxIvZpT5lAHLTZJHex6kDQVPZqmqng7JPVCpOW0bbn0kA3LSpUmh3SfZ5Hwoq1b4HI5Wn8
TlC/yGRseCB43gKTrpn4Qm/DAb4mUjJOTtZ5M1tXQ7HcVg0W65HLE3fkeJU048ck/9l9V/Rzr4jF
UkhtLGBRuL88pQ1Y8hZP0Lw7i0QcQVVgK+/ygVjybSIhlvE6VgLl4Q7PBAWSOE8iaaSdW0o42FUV
zax4lRzRijQa2pn/tTPBZaKjjnSH1gKa4yr1rGzCLkgMPs/Mejmv9fCXM9Km4v/qgwNJmc8+w101
vzAkS5Q8c0RtRF3kHNh6vkgZanMxUTyospECIdREmIXK9fr4FDWqZZ3nTIlgm9JwsvmoSz/Q3kit
h80ysUXkFXfoIqh+9FNsRgpqIYgQsSC9AzXvIsRwXqSbmuH8SpVr7B5Ipk4D31QZCJB6CGeqPu9f
yeKj0pOIw2ow5/+PmEUXdWPS/TtaQJCe1kkRzYqw1NEbC79B5phyIRDyq7rxfpr1jUGG8uv1rY17
ZjYrR6a/ueG+X/zQFBqpFHE2tchHT34mjwthTy27p412iEgH6DwPUJKJNaJp+88fn6wRpIMiYf20
E4OpaU9Eg8KbDTQy/ROWxnLyc+5McHlL2FA9x8msbqVJ7wbGE0k91IM4N3im4R0BX75GnGSIc4Bo
Q4aBwa/IC+MmE12zP1mYSMR15n8QGUKg14rY5ve5hYNS9oCt/VVbXPiozWv2nmKQy96uMrQoQdkj
njlrgKQCtLDrbEzCTbJmZ/RJcbIEiuAKi3+QVgy0ssTJ2CrJSfoBonlZrjyt0bd9DvatXvNcrTAR
S2vy9ZB2NC2Y2Zur7D8DRGCUB1OXBjDZU0GGkHxo0dHrHOdtJ6d2hpkxsZrmVIvItXuaAsAytdR0
Xzx4rW2xRrfZbibkGFAaUlXl0F3+GaNPHxAlzOux1nVus7GdvePZfajHKHxc6RxEKLYDp3atUv8k
QWmbQqcTv4PfV+OUf3mjyXa/86rHdlB7vbHgI59orIKR3kVdABNhiG6Flrbne+s8nqfASG2V5Vvy
w50Dp4bT1FTFp5eK/n0yoqFM5IIpXvu4rpQw4YjGpXFBygiTA822Pt5G5BHZDMa6DCvfzAYByfYW
bThTUyouZOxqsEexTg10MtMCf/riDrXIBdf52pseresNW4Yjt+dggtH1jMhr8KjkNyYHJj9GDTiH
6B1l/2wJ/tc2/p5sxFLDfNJeFJ8HHNCgzV7weaiFqvKQkZZ5eGt84gi5ZCq0oYQ+s5a8VtWA+1cs
dGQ29zhlbtMzBu5c6JxoMaqxsEL0ztTKm8nfd43UposIlbKXz65rHjKDBkEYQZ9d5nboRMeYkyUK
ElGKBHvnEYB8rK1BcrbDX80j0dhQV0ec2E+7UL+AiYJlatm6LmajGZd+uWjwBoZbbo5lqnsZWSxL
R7eovh1uYC4RMwdTjiroP2oNU1wyh8OM80tHbqdEH89zs1t5PXMZBIpsgP+ybcg/6Km4HX5xDuKw
htGOkoIZ6Ta2NpMSOMxqzJwAg2wSQgTRiKhe4RNE7QaCdDs7DZmvpfVRp1QWRxVmbu2iWdAU0FV/
FIoPP2983gXxj6HgGAsSVh7X/2EtoA3/YSyz1PA7q9SyTJf+geyaxFeAe3aczN8V+qxLhAPcggvx
rdXJDHZ3L9XN+erwDvQCinlRQf7mVq3fXSHacGr9bJU0MDqanez3sHz8pfIpLJh4P7TlXnmKHyqj
gEi1VZ+o0TWcEDbWrb3ZZg9LpO8g466N3uhINtMzAsN9xOMeQYc0XIb+zRCiuWThSD8k4AJfYdam
ZN2Kp/tgqLN0dOxw/Tdw5FvGKBczOYQAmdJBxAALYHJQly+4VrtwN/RxVc0Y0ET4h/vLsVOSrVEN
XJojWOodljaiiQy3L4K7mtqTSrizfg+k175wGM/bEUIE2qJWvbDecGeu1bjk91yp6llQICc77uGh
BOIbigdL8YMkJv7/qNWnRLPK6topLRjfLBhTckzLJuYStD0NNoqtJBBEGCP2uCPiWm4jhcAsiCIQ
s90A6EYfRqnWTv0xWJh0mciIdJWYktnfXGbhDFavOQJ0Pmab9oH1vWPpANWbinUMtKoDtCI9iVru
U+M9uvUt+Dt8EpktZDJhxUhkmDYy6OMWY/Ax6sAsqbcfmTXBtHKPTxOcLfrj/8pmbYalBRoSvjjN
fOCDs8b7TTHH7Jxy1yWUK0pCH9MAFbXtNq9ujMXu7QrjnnuyrsWP05uXZykw/PVmSabLBXoxAw6K
9gAMNnQSwjbzOhMa60B7WY8qBAPY3hLRXlDWUhB3CrBXsLW/GFnjSEhggFqPqTdPzLZrXL5Ajo8r
EkziqRA0l+sko76MC5ULkOAyXgFPfql0OfmIZH6PllujpOWT+MubcReFw+4oKPhhrAMVdQy5MLdu
brlc7CEKT27etx+jyh8oZBHuE+8q43EKjfwuDcArdt5WGZkMSYT9SB8WuYroBVMvBny1lUpcrFvb
7X/+he6UFKILdnAiGwHgxpFq8mi800upl8cQjs6BYIbeoT3iSXhUaKQ5oyuxKdx0QuLvsra7TgPF
Sk2uk1DiYq8nBZuTDwwWyRCeXlgSa0H6pPr1bG+2jL/bqutHMU6ol26thmBaNLJ1f55QMgsAJykb
mbrq9Ab/hXfOSzCa01VHgDwesrChkcUSWIeGJAwhIFbHFWjlR6koxJxrMgX3QRGQC/Dk4gNI6w80
7H9/Rzhpq5ht2VyNHRxhcjkk6NxRRUUSC18sphqa1UD4FqeLNh0bOk+ORqdphP1jwvcsx633JPiZ
Wrvxo5Vg/CKZ82IsL3dyBbonFJPKLtfHK6G67UtdLHJ0qSpZGg7+p+7wwIvQhlQj67NlxzCYaUsZ
4Yec1X2Zsdzcr3K+RhWnWFqDNVoAMkxazEX+HQFMrPAzPO5+yh0dHBDjHjZsRgODDDafVCTp6y5g
kWfBCH9tPRI9LosLlyoc5H4goXliGKewzMLiULwzc5GjeA5Ib/HNwq7Tc+3X+XymIwIkyTPzfuIm
d9iCympCy1+TcnXRF46XqT4ckww2uOllPB4mcEIFw9GPthScMWbGjmaiZQoHRH2/IfD/kTOX0++S
F4kP3jkrjP/VkFfpwyJdulOTQo49cZXkvwIEzfihIVmZut1Y8KS39fuVhuKwB9ck7YDXb0BwEPJI
p5q9a4W8kHIOVfXKB5EWMO4w7zVDjfRV9kVNPSlv8H5OOoGvOSh64/Ut0EbFttTQOYATSehriJFf
KBHMnjh57SugWjlkF6JsAlw1TBtwPrl/NTULtemVI3vB0/GTC235Kvg38H/Q7eF6nx9UvVlRq/AK
p7yPe+l7z08N0b4dceLylM1N6DNzqDNzSk/qKjZ6Quqm+GywL7QLhh0UTgFp0LtFjYJgB43ks6c1
5i0QcTr6y9kJXG1n1Y9N56DD8NOqbA6JWbCByDaO5ry3ucL4vkUtamLRczbYqy9qUIffdFXuQ+Ep
8EA/ct6jmXhK1XiJdpnyLnftCqVJqjb4MAmSrWokejcOy+PjUDXXJwVlX43YvBmueesAPK9uLNts
zjlQ/svwYL25HOzdPtlFXXFlqbd/LczXdDtY8iOvGOlyrIX50ogUf3bYJZPLhuusoySL2A/7+tjw
JPSuRO0QN/nRYB1PhyLXgQzBeaT0ouZ1MN4uSVYijZoljtStDX58lq84Sq9pfLZQdVX0QvBVb1SI
LEzZ/G+K7gpQu8TZst5F9zFu28uWIotlj8K46h4MJtSj9uUeN5yoqKEcMimKwI3WhrLIOsm6RFV7
aAv7IohwFX/BxK2itlvggRwm7Jgi3g0ycbHOeaRsjc0F/kVEYBl2yT49jxHJswTlsyIJLPlxnAsM
/FGWmu1IOb80az5F5FEpsqDhteJN3gAzt9/LnJRlt/QVsj4GAk2vPO7crsy1nSm0tTD56YPFZXqx
WGtjh2lGL2HxoTyyRGHCudDRLsdG7wDfmnWKsnAqKqX6YCovJy4KA6Lek6P8iuCx2G6dWi7k69xl
qMZhTO2RXbAPYrsTQlCzbwXHx7on+oBSgkSLp5asiZPr0r6/M2JQsQPnuz9IepgRv+YhdbkWGtvT
c1ot7X1XmrLde81vYHqZYgLi0roaSZ26nsY4sjUjntZXDjTnTly/ghU5dY/Rz2a3spSYiBEA7jzN
Xi4GmoX5+Kl8JvtfHNILgiuucw5r11gvg6Ee7vJgDnYD+1erVOFRE2TPr+u05BE1bEKiZN1StbAe
fF0ZMWOOHNHMV7siFcCSP5/YHGB+IZK1iKDACLCv9Vb2AYngAn+oXe41uYk3O1mR6ZH9J0CI8T8T
3vl4sJ3fkfi8taaUtVuk9WTCQReGMDEYWVK/fah2znGdamtS7EKddMg0C+pPySU6qDiIWeeoI51y
UuSkhuJk9D1NO4TV/Nh5mOcLYKAJboqygVgO9k9Ix4gbr9rFgKTOVqTAl4mn1UF/jyoBlq1ORGdy
gZanQG/0QdMM3WJS825mIcvRzMIX8AZ69sIrtmG54ECWZzNFkXNaAfNA9PKbqraFogCOEf+vPKVt
+3CYQpUhEJeYLhYxRSZ3YCuX3OuK+tAXu9ZJiN1q7eE0vco1m0JYk3+9mWtCTf1Kij3tWdHUn4Tr
28LbeNF0kaNHbnRFPib9CDNcgZLMHmVHDiaGno55mO49A5XwYj0XNJiOXZ/PeZv3+2BqLm1Q2xLp
JQbBzv1RNBLirbyoipeBJ9O0VC38WXps8E1kG3QGYDa8zcAP/3Vl/DLUdz9eylwDMz6O0bR1klku
rmC/pPlZGGxcI3Odt8yhryCD/hIJ0qO0clZ/7K4FDJku13eAZnh7ZGjw47xbDfJUCX1dTQL6qtGw
SkcafIEFwV2uAXPqCnWpydzdrN+4ymOrvE0DelUE28iLpzDnZHkYpXfi88liV2wWlidiS0PlIgQL
T1NoqOT74L8y/MKceHKOOF5TUVagy/Xz5BL9nlqBD61hPSVwz4SFLrKJPnseeV4wGmHkPX//RmFC
2jRUZcA5clBw5fqW7ZtMp6Gq8N9CaaDCYcLnuS3nCYVDTTJjLuocP0DA0ziRvdNOd3tKYI1kkhhz
3DWLZlAEoDXZmReo/xxjq8o2Z5ydj34E1KHdJam1SbH+PBZH9Dprrj/rNpRAc6fhljVXWn0vMADj
RaWDzumIETN8dTAwH3imN1sT6mXrLQOAz1N200bGJhIyJ67ZizuueyswTXyOzdBAFuk4Q/UpM2oX
bXjb3s6B1AVmnp9uuwDPEkEpbNbelfnUk13iUY7kGWwQP3+W8DO52wjY4JjfxO94YowblvZmYyd1
+iOKzP9OPAjw6TmYk/5M9AXVvx6eyc1PPjc9p+3Dp6pTPMVKRObiY71raGgv4MR15q476WtLfpcL
hLbhvaQwxP3hatRcbC8n9OpyOsuq02NhENZZnFFG4eaMaQBGQr1xZSIsI8TEXYCjqt7mUK0uU6NA
lJRtGnUIF3rmosafsF/hGfvttVhXJ+07edC0U9+zvdTbjBmJGq9ybQoCFoZx90OnxUqU1KvDRgpa
01VWyhuiH+4kd966QrC8oU8ITJS7bAj9dT5CP6/f5UrE/FzstSEA4gGbnAvL2On7qPEdfKUI1vlq
wIoj+Gf/zJRQ5RXrVaUCGcHbIMCGcsbcFjUXZYnqqk1n+USwMsUIzmTg4flVMKvBcBUqJoqkbjMr
sl/13O5TzDGzcaevgeIQH7C9AmQTJwORazWxuHDcPPaIjd40hPf0rkRzO7GK1LCyPR/jf0WBTDpz
hVrpvjEmAxONbZli+VOdtU8vP7RSTSbquTrBotGiKVQ64PA/VDG5f0szj3/wKPRUhNCRyS+hF9Ws
PEwhnb+lkekEgOb3LngTqRYBRE2rF6a3VZ4ievs4P1046C2+uEvboOh96yJdXYF0toCiMhbdi8m1
Vfy6kmmmdZAuiL9ySXwY0jXZjrNYe1XXvp4Mah7lMIFa2+00smk0P6yjOUQ2yZfXxnml5ehdXY6r
C0z8qMq7WAGyYfjrTHSE1mLqSaES9Xlfl5+8YtBIAyvi29ZBFbbnK0rgN4tdqiBT1B6xaUl94V+8
3VYk1/w5p/SSql83pLVEqiHrPsnLmwyD3IxgpYUFVHD14oGUMtL9SfkIuefVqSM5bkYR7+icEQLs
ieQBuUUsDo2HbUr37X3IFgWgWG1us1O4sef/pJpB+2OXl7Vr8DyLQXWexCdPBFioKAgi+Uk2HLP+
wwfcafXPYxw9/fCqxPCcaR6+epc0mEtwysHclw0oCZxgcRVHbzTGOwT9nWGvc+AqAc+M7xx82lIr
0ItxOt6EOlE5Ic6rUDAN8OHm7IkSCy9xCXIamGlGfqiJBfflvEmPDRLh554ozk+0O9msbhjuEJ+N
+U5ks7zOvPomKTbsGQyJcSul2gRlnsHrBNfo3eslxxBtrWGG1fxJ3+rOcyTa8DmV6Bw/FOmU4p9r
FoshKzYnQPUrlW5+gaEOe85gGGdTL+ylNjLIccQG2i4/ZODO2LwwxrBzZIEWJvj6cnTM4ftAMgKA
oxuwYYmspAQnF+nbel9922QsA/g/yQ2d0Zzo+iwdfSC7+4Mq/Tpht0SynZXdUjmwY2v1wZt7Lxn1
xcYGYcxOyxNpPlECPnsa0dk8VAWGf+tB0clbnekLWJCJsDrFCf6gR8Xa619jW7OODuNuAFBGBJh0
9mUL6weDc1LYiy6OcrFuUMPs1fFWbxBE5inYl0rnnFKpOtgDxH0/AE+5sarMZIfua0zhcjl2h3ng
FsV9yi6BRHbs6vLwAUSDWKMw9iTMBwXYu443GfMGPzSMsoWRvKGTVoMdN1vZqRE8yMi4Bs8+bjxv
BE3cQhq/qSPHcxs4nQzsaJI5OmuWfSdzLyTuLQdZxP10d+cOLhA4+aRAvBeIDfXkk029EMQjheS2
2+IWUoqEPEQLNhxjk//I8Fw8iM4BSge/H8HXM0JoeW8q792kPm5HEHh1qeMpQCe/1eTFqzpr4hAE
vhuPOcR3dcpbqUArvl5j8JgpW7M/TJaGxFxITR7lQ6zUAm1Z+NIHeO3r/+EWg6M84nZh2QWc4APq
JzbVEhFy8SwW51jtYRutgheITOvrlMrwOwfZFLdjeNIaEmDyjw6SIkNzDfFuyc4CzpTeOEPKkXqy
XcpG+nkX0tEIUq4E7VYDqMAFcuZMIycXbLBK/1wMkvufZrFBLwvqu2MRA7f+KVyIatXp73rD82j3
IXmAzaA/He0H0WAmuCc9RMVd1PGXGeDVkXVXazT/yhDttVxbhDMKI9MaBQVuE04/xoYwrZR6Zi+P
r/DznWLBWz/KXfC0lmiEwQIr0ImNrXC4MSTsSu6DosD3387XBAYfKlF5NqAQxrl9SdiKblbmhYm6
0EoFLomjvknalgXkxd7ro5HGsnRgkssPng+Z9gDAN5lCUUwtTNH7VyT8mnRKYz5Qr7+kOnVq2uEP
uVZUA+cU+sV5rhdcZoDlzbhMVBsF5Fd+dNtE4l8Jhq60vBXNpusrq+Bcc3/qLjgm1EQMKGDBuAPZ
uz4yWAM/4/5gJioHmcXHkjHAOelA0ACjKRzf0kD/M42FYaXvRemVgL0RX88FHu7AgCTidH1wbXzK
VXBgt8amXr/R4FZkQHEiww5kxyFDKwUK3u50zX9TtYhCtb3/OKzmvgHrBgJ9e+KLamDu5sjufweC
eaHlz5zSFMEthTcwiKmNyrBzs+JeLaM8J4ltfIBuY6CIv0AwxaNbYBrW8OyyQTpqv1XJltfzCo5D
aCx8CurZQQ/bGwaM9ofi8Qwnh6l19e3dNa8xAscqOAXitNPKFezvqTgfruiB9hxH8zMkBBIHmRp7
hm+Q+VNH6QvCHaSK3ZEHA1zjnYkMhOEMGYhZrG6rYPkMHdvaE71TdKTTtSeljKDoden0c2m4GiET
16wuQWDvYixDGzRYP3N23C+nlpjvwSXaQnEnbt5MCeELrrQ22/LjcQ6aTVVy1p/vI1su2evtT8VC
KZ4dAJcFLVriW1Cx3636wkR7KfEma81Sa76M67KgM676LE/VO51jZJyoTvq7W7EpMDGL1FiS6KvT
922fqhyQ9RscDrkhmMCMhbqBXuaH08Pl6/brk9KgPt7jMYQGiNz7g63AU5vA9Pr6W8wW/bsMO9K3
pjfYvB3ln9igTfqfXXvqerDQA9NSWjE4S1r2tvFkSes+4ktnF+fUyHkYcCGHZWH+XPs+lgecK40S
z2hqmaZvx4c0zt24ZDqwmXdpHMf3mLiUv8Emgow9US2bW4eo5l9frLVhMM+rhmYW2exg4s3URfoI
JniYH4jlF7FbZ9r4OA04Qfi80Y1DsisxOk8EncknDM9MmH4LNlYCEw+CPeyyrVE61ZB5mE36IhzP
Btb9fzmty3BK4ew8GyrJLTQai7M8TOgWBGoJtB8zAwOxpFjYxAIf6N/9yVE6a+xcLmcrxO0PQf4G
WyHj8kVPLD1/sfftu7/851KXh13UG0cIx+lv8za9QG2byayhQxokRJqE+mm/frdab0Ng2v7Y4wdd
ASJL8xY6z6rZSQP8ufqtHC90Rlj1ktnoSji+kxRMHNn00kxrJM9byU9L4KITudLdgvdhi/C6TIjf
KcodZSrAOWrv0k6XTBrh6V2mJs4KjuSBgpEJ2tJf1BoiAZsgjXWtx9mbVoMjp2SzsV9k9i8QfgdN
I2zJZ2bXZamNTEBDvxLu9L5PBWeZobdgETphooL0lFsObD7NomCFECyv1TH+lB1Fn1K5fgJV0WuI
iPZ9BD5sz9kmlH6JHZM/rNTejrf2iQZ5dX7yLm7JX1NDCKb7CYc4xWFMCzIIpcAV17uNG3M1wuNW
ZWskcVzLhkNLWMMYLIJh+fQswwj2elEKhAY4dwSl8Dz449R2Pmm8sZphz50R42t2LD5o8QVaBaaH
8DJRgV7DToWD6gjrw3F3kH6ihs7uM394/GEgyf+agX6D34Zy+80Ws6ie6TRuU1VQcuhZazLdyYm6
/6L5TDCol+xFcTkoonzkgwkKXN88WhbTj9fQ9lBrzgqZYhr6yZA85zM0v/hrz7jCYE1r2VNz0sc+
hKyjp7yR7M51/ZXb1Re/UbsBAdTCoT/SEiK65ApOz9ktT6prCcYewy8g701e6sNLm/bFQ15rFSgt
eEluhX+rjznB0kh3Ia+kkO4lVD1pj0bsI1GQeXdxIWIO2zdWuv/EjjPfH4T+/qq7FcVrdCxtEpdw
2oITN9fIPve3U8YaV8ZxRG7b/aVxROw9HjNq+3aEA3gXIQ8lsm/V7MSKQ6PD5Ce51tWX4vW0yoYy
LG6qBAyx16W9VDQaLxfpgxJ140Iy0ZuNuXa9s2jfQ2i2dq66b6LPkgu6pCRviYoVmWNfNhP0KPDE
fKwEyzLSPfo9PbNq1s8ekkpkCnTSpkTR750BqReMrmpMP+wLOHQTroWzIVgcafNZ7+Uup0IVHqDr
Tp1kWiaS077Twp9gtk+euI9G0iV3S6MyRK0MjdvHyy+xaGteUdvf00ZltPh8hTwLKpvMMJdXGEan
6QZlBUc9wLFMrx2HgjCKevp16SoCG5AHbvdXooND8jol2+I3BWBBBL0/RfIrBuMGaq8UVtF06ZiF
M0m3lcbsWpi1GkB4e6QViONvRePnX67HiFTGKX89RwRinsHtz3yA63UADGfP2ePlVfmQcwrxlndX
0of5fJ3XDDQs91gBP+N0sBESvLwQUEwxxRiBxIx3OC24g1pTwnpcjwjsv1KlNrVVjFG+Cik+m0Of
oqnJExGVWCB4V0dRLKJqHmuzD37TeXyVEEMQePssNG7zEG5lGaO4zBnL/u4VYJI3XdXvM//6XlfI
eO6IVLqyufMSjD7tPCaoV1GsQZ4MH3zmzTvEPy/J/ZVrfe/RaKGWbRegI7mVf07+0SGuw5rvXyCu
Sdadx0P26jKZQNfmQ+V9ndQHJh3i7GdTbEDxl5+/8xxTooOeuF1DQGbqljYSM0tJxvAJ8YZhqx9V
++1HJ8diJyPCefHduJ5HpUL1cEUiTxrVtwV+h7Qx42TKYFz4hIBx5/xnpHVOQDSET2OGMDFKFMuL
GRilI98NVarlaDYYpTaA51N9MVeV1bNLYn8DqotnNSFas7zL4K5JZkhifnQbkeU1Kxvl+Shi8ikx
EfVQ5DZ3XjBjAVTs1U60eXohw3EQz/6/jMz5oU2QRrz5T1Lo8KpOWhyQA6SGDUyxJGOS2JD0EU4G
kQA9ieBYuGOK5WLaECK9kprNJ6JxfDqoZfZ/hMdAXm61PY7cb4Wti/IbMVTUr61y87/2EFzBfNQf
CFPGJ6WVGQ2xMfFw/MsPd7pOOHtRwsU1XhnJTXnqxZvnmSuFffZFNNL+Wj9EAXU3YZyWscNvmiP4
S7Ycdm05W7JsTK/QtbtVR4UEb1wIjNqYIyW5A9OXtr+pvYmHf5y8PDNmhePYWEWI1TX2V1BesSNd
Un8n1HfFp9MyoHTld29soWerUXo71SUaJjpxCJEQ+RxLDzMcu3mvwFN8/paiRogAG+uFppul01mi
8YT6uGmxL5HzRo6XEnLGbRXbObsZ57nOpOSMX9vRiHR2hFwfx8nTDx2XDVpouRzvRoqOFV85Xfy3
xA2tgaGeu7W8T15MvaTD3jjGFt1xTpWPz2Yo1hDACma3AOamuFz9cIWA+BG2npefbnk9+xYjRbcz
jHOTw3/4oRt4u38QmnvYcC2ZHcYQhyL9ux/8haQ+T31B+MNVIHvCN8PtyVg+vZ+NgchXA+SA16Yv
TDaofTzzIDJX7uN9cI4UlCbIZHQ6cP985rFCvtL21vLrbCYGmwXBupcQjQozfemih14wslqghfVB
NuGxjoWBDuWIAEy8283KBvAdD76WcWJbwepuOWljbAgiuG5Kmg1ASP5YGr3WOs9Zi240y4Gh2M4q
kRh+TsrI/FBG6X/wJPHoAv9N5tsu2VH2nlYgYBPVivjCVXyTTwmg0g2okf0qhb6h78fxjxM91Wfs
jEQRz+sXRUUE3s0EzTQARgjr7tjQWhotQnWZWJFitJR0LVvwZwYz+pT9D4yrB8IPm3oLZQzl2+Af
p4c2qVwQcCVBoFk0uhkUUSNE8M5q9HAiB72DYHidUWvqFAGLZNKcP+fF9Ur8FykqCmq/f+W4Hn/w
F3CDhIiGBbXYhYYtWeE18V4VFiojCnFr8aF+kTePwUDG82S33dIH+KHNMf8B5w1/8n95X+zI21B4
BEjialwwSzG/T1xHuOFqQAbTyEE6P2oThiRvOCupV7R0AXhI4K4quXP6CndRjmDxl0+V9mZhx+NX
1cSbZZWpDI2lusqDZjCL1+mLEfpn59Czc8FzTUtIxU6SuqDy0t7VNrshpDKjfiZkVbeZOrDgb1w9
PXeLsZIaphWO2Yj4FTVhBNnxCIeFDuX5N3FlOeW7lpKpntvwY6vRuTM3Jas8Zt9b7flts2KutvX0
PGEN049HV+GGvuohUkY8YnKFpb0g0krypbnUPhHsZL+7Hd07duyJ8HzizAAZ1gG2ZqFAJETkY2Z/
UqckyO9rFauAUuVv5dPZ/arAV0kbUNqR4CSU5ee9bGkQENG3r/v0/c4LYU5CP/yKanNEjouCIzeu
a60+faPmS9WqgXaoTw8fHAO/a6pBsQ2aa1Q1JpzZpxk97rkQiF9o0BjQdCyYvvbsUK9vIFF95xzh
CvtWC0fmqeP9Lx5Lnjh9ODrn+GFs7Sh5uqDj3uT3UycEpKQZTZRXnk8Ukeo6vgxNoXhfJ3JT9zyN
mfpa1/yimUM7fW+IMxLn+OtMdQeYs9HgbdvW++bZ8swgmW/FCRkX70+3EpXHBL3BuGNziokaB6uh
YooQZfmwq4C5nN1ka2fEeMNP1xuohPaXQzdnhO8wEMkzlNfypZ2r7zPlcz1KXQymOLnjOfIqxEPb
HcQXf9dB8VbXMLv+t0+4hQpjowMM7zS/bgE97wzS4TLENtgepfXjSnDhooUYnLvLZFgSrAQD8sev
3PHeR7LzAV1BB6oktF+U491A1cTh0xxc2Ja0MmHLs8DQj7fFz4OE+aBpXSQlumDrFBFpp9jsobV/
tS/vJse43u/rqnPldOoqQEcC33YGCk7EXU9AG4yKIWKuq8C9dpOEfSOg5fsh49bJGbAXwM+4qISe
I+g9G25UYHsA2ulKGFow7qGFDnyK3VsDUSoTj0A45jGckuIQptXVuywDKzviyxSAiJghe4pEAx75
QpNzWITsY31Aowf+rVCqjeBzwaZuLH652zzy0piGFzwh02YCMo7nv9KTXhjrXLbwZpL74VI1OU6x
4SFKm4vaCvGEjvnqoxIzkUJVz/ZKLKgeeMb7YrRRcsowqRWsOCgZ4LzgKGBsVv/zOa8kU7/ps/N/
pZuMQoEwvc/AhRcplm3QG4rn+b7HNN1p7I8gNHgvzDO4TlDTetkBBLXykR9/RR99FIj5+ExIaUm0
4pa10pleg9OpD9+B1JeEwEF0Hk9JjaV/NB6ykdWg0v++nX3HlndsK9uXyAmGYqdRsLU66dPZCEBN
GfmqJS05RusVdzeBgxzRMi/9MdFopVF8G64FTVmoOI83idd9WPlyt1Budm7d2m2zFid5tKH4dtn1
GLboWTWO1mWFZ881p7oMoF0KNt5OndhkAI8etEBzlhlwYkMmIIA8nb/RuwE72kvZbmldYJWJOIZA
k2DLaDHtd6uQrn+DV1edwDfp7DCPE0sLD7WbHNjno0su6Ld7MTGF/EUT9/avWqFD9jJcat+9smFy
UeKjjYIP4eE/BwW7+EMUnNQIUrhI1sxyUhS3x/l2rgh4HrZDDRjlze2qHE5p+YcDB4E5s9YuWtOm
Lfwsajfqx4ut0JT9P5EqwfUB9pc1GUNq0i87RBHN2NTudb9cfYefD/puvXquqQlu1QQUNdNRrqxO
rFW+BJMFdjyBNxtC52hOicDvpWjznBKqAP1Z14ddZa/iqxTF4t/IaAWNE9blVx/1B5OMkQcPew2N
SGNsU8sbiQysG9jFrV2nRh61U5O4qbeDtb8fYkogOzFFjc8PXc/16UQaKktd8SSpFRQLhmRq0o01
rH5jo8D1QdNCOPkpuaUTTzWhpCZL0GxfOXhHqW0kRq517suBZfm1CSohWh+FEgPRfx1WVqePlAyr
Za4AVhc0BcXrqnyKc08xYhP0D0ymznfg0XZ1UhFAsskW/bkICQxZ1LT5WwotgtwEzmvoqNY64mNk
EaIqY14pjFmcA3JlNNw9S3qr3Ko7fF5J7ZC8z+scpr4OxBOffMOKoS9jJjxoA/Aiv+naXGFPD1xS
D6nbkQPFweJXXKd07SEjekes6O+OvXIJ/sLzBXr8emi4umD7UTL2SbwkAyeel3XmRBvYAmM9GQh0
Y22b9bLjHjNtuoyaCgMblMbQgFhMQjXXaOcMkX7Tn65b3oVaLiZMPowPAcHWhA0zKo9Twiyxamws
QNoJVaRptN137htaN4SCppxEbX68FAxvODKY6FK8Sc7f4aILMLrVaKKtO8XQR9GbBpSObiCYiDhy
1FNuzrPGyFVZ/V5XXR4d+cocVVBn125oL9VuNx4R01kOXPVySmVRg6ScNgKMDhiD6AiLpIq+ksSt
NEwAZnXFJbMbVw4oynyYymKcGGqJy0EibuoHnlxE2F8laNCcDsTUjHko9Yy/gY5nqe4B+Yv8z1nh
xNcx4qNtmTonh8p+WIkGxxdwYVxXeSlYxOv/ia+3BpWHrOlXUTt+ZJZ9JXwM6tTnx0kTHHLvLoeR
GuZUKhQ55aR6UdcgDPKNi4ePtY2UDxU9lwVlgOHHqXquaoIisy5cZUrlqA6XY5GnAQ4gW4EAnhnF
fACSkdBjxEa5hRA9Qd00KRaTezENX97x6w60EDX+sShwptZ+vrVo33uF9vu4GmhZFqqPafSfN5Nj
1kyStvfnqZvIJRZMt1t9EX4Tf0N1jaNuJlIZu/ZaH3b+CIACiMXNBH9Ny6YR5KtP9zMxMGvemnhb
ov8B7Y/yk8iVEgeTHHf/8HWvDAC061zAtMEcKoz9pbulgIAhzs6Mxo/DIQvuDpS/1029/tBb6Q7R
Kb0Bvawfn1liKp8uMYya8XRSCOot9OO1vAJo63e1B/cI3Th9LISBYN5mZ4D47yVZx3M89etcQeLS
/3Mcl4lh/8lpXw41o8nzPyDHgiv2Haj0MDqSQ/qv73A9XZYwT7MqgNHjXE/pWW1BkFlqpeNyUd1q
CeHSMZ9n02Y05TToL6HPO7z27Y/4aXO/7u1Hq2kpdVB9zTsL09s8ypJsfEUge1fo/NYFmQVeMzDN
gOaT+pgpTGCsLzn1VB2TKtd2wqyW+W22RJYjZWkC4keuqID8uYf/hxdj4jkiQocKmae9JS9hiiZN
4eNLOSZDTi50wJgJLCfGTHYXTziTXAGqXJBiTdi2E+hKU5PysXSIWC1uqkab4gQbk192xlR1bNIo
vx5ngRIDNCf8dEsuP3dnXGN6GTOOUOZHA17/yUMm3LOXq7oZPtBtfVUmTZySAFeEHEXdOxZhHzPf
YBCCzlXWt5MJ+vEPtn7OuBQzykL/6Jt6qp9fvHcxgwReDeituN5ztnsRVRIrWLqIk4Cp1AWwFfvP
s60s05BPBUirbmgKAmBy4bGUE5rYNlhDQe0Tu5qiWU+DMR4wAj15hC7/jGA0Owxps+qheEmjV2X7
TD0avaCuphV7gSwzKqxJMZx6akEcp7+HW7FlXvh5dJ2pSOssHWQDfHr3M5dJ95g1WXjOF38gqTFH
Lq693QBStNpOd0Jg2wtnA87n8dxKfJqUElJDieflYwsoUM0ywu2eyXeUU2wpMsnaGhu8Kt9Tk9ry
S1uKP4fYqMbHnnat9AFeWmGWQ76nA6vW+YKeguRPVEMPegiiQBufYL8myZg4AbArrL5ObtkhcpIy
uwW6QumRt0OzT92GJNWxQar6hd1NN8h45lstqtjcM/r6iIsvJjNIZFNXG3w1GRppPe3M/Jcos7CL
gbDChLbWnoCl7n79Y7k3zceBk9hWc1kYKgRtOeoENYkvEiY0u6zJLLvAOey6amW5z2s8dxvCGxMx
V3y/6cYnSAA5Bn2eMe9AHDfq/HSwWEK0pwrT9zNSTyzBcULG7jguIFrUwKZAf3PyOXPsoVWb/ejK
4smYXhDO5tWYpwRi+WmhXNSaIs/MNuwEghP5DBDEJzhMwyisRE23TNm0zY8yLf+J9IrkbHpGN/sT
jK4l1ZZ2kcw7Zv/Ki1cQwZIPt3XTmKgfkYrBIyQfZODtuPsIg4HkTZRFNKr8BPc3sAEJpPDdxRB5
szUIPSObRb75kFXCc1p8AbtnI6WQ6ECtUgSvvmmyAT150PtZJaq6XQgPn14Hc+4pmLEfMouGQYgF
4EMDw/I1tT4tEr/cESOakGNI3frLKmYlIUwPavlLjbOnUdmo9prc58cc/gMa/v/rZtWci3YWG2RL
azXFIXvZg2E3j9vIudOogPDSHznRjZdW6lgT3N3ol5618Y3GERXUu67YOkr2QIh+DRxkAggE0jh7
lgxIZaedDvLtIyUMDUioX4xBRaqafl/QHyYlXTD+IK0CM6x4zV1hCltty82CpBedyQt9CUzKcjVm
URScILSHnqhQ3mN9YJrobkx9IuwNHUiuREf7fbRwbf3yMG91VqdZ1L+g6THqeLcFxxbOOpB9BCKf
/X79BK92OMpvPH3lU30WR6ShytXkqV34Vnkr/egcW9Yrwo6UW9hQZlTsLStiO4Zl+Gk+pwETJu01
eS9DEaI/SCtWPfaTtygZOMab0QTeuGkye6L9QUtDljmoq4LDPkLkADWPvgk+GX2sfn/6p+w7ZtPr
G96f4vtErF5mfY4IG743hzLwGekGO/G8UlzNMssAet7Z19wslc0FEsC6rAQy9p+IoUrfVsgXrwoI
wLvVtE2w8BPI9Sy93uypwnTXfxYKu1QcW7Pjjz0dW25OxM+Gr4tc8FVrbRWfmDG5Iior4GoDqt3t
kbq02FqxRTDn7owsRZZZX5sneHnYGPKEEHad7CaaNk97PVOUf7JzOvPTS7iSJoHDlU7DtLAFwCvR
7ApRyXOzv6Xi9MbCINeAq4ygy551LBW3BPwdbuOAZ+IKbY2fCL0J1n1NpdIjRqlcw5LsbQbaT/fY
yD2cvwHsJeU/A6bfa9cztSX7pdgsdTJHI/YPXYZeAd3BgMj2/vqRI+RsjjVNWf+n0v01Z64I/YAj
wmhKP3ahhe/bBpcEdAnr43KIIz7huz1yDklPehd8/3Xin+d0YnjIS7ObHbUDkZanOVezLOnE40yk
rt25eNiogJ06ZxY1PiOZIxUqlHxk/4TDi2j5SnWaDC2EH31mWS5mKUPt9NOWT9I40qEkRcG2KcGi
ltE1H7AxQ+7sRk9G0RN6qeYNosJ7yZODwBgpDW9X0SjeTnf5zZf0EG+dziIbia1mS+x7euyCI4Cn
Brb74CgiI8dOcY6rbRJgCQRypt5qORalp6jFeSVXfMmN0fLg5ZP3drXsTkQ+Z8//durg+P3qW1AM
yBzWX4yhGBkDLTajPt6VsDv+Pn/IFB2TgbyUwdRpH3A23Xi8t5EhINvZkZ7EK1ab82grD4UMb2US
48LbozTo7qZgoeB+4XqwkYIhPRozlvl6HQTMZAWFNHm7ZCeEbdtjAwHtBrP9BWLJh5IXNiRNTwM+
FtwHrJf/AJYOuNBbJaG60HQsHXbwQ05d1Tf7VJ8cebt1Q1BZm3tBz4pGqcv87YSpSC2W8h1kpXeb
0E3pE67Gheuer6feuWbL1hzgI+MkhRyGka/r0RJ+zKHxRbwZnTdkug3Qby9hrTsJGPWSibcereXn
E2DjBtgk081SY1Pk9/su0v6i2tiN9LjXdWEMmakwXDd5ieOGezV7Z26f99k9+2GZDWJp3mRxh+TG
5vtBG+B3wUA/17xWu702kTp8TEdD0xp8bUwWhhJHowO1tkIKlNT8q2Lc+DnI4/8o1pe5s9JLELrO
TMNc537XtgWVYzycQJq/WU4juEOsSTf6lBm1SE6OeQedyZEFxBTP7kw6qCIVBsIII9guPbkxIr6t
9sYOfv8FRZApQmeZDBJY4nDDDq2FljcPvcKvqPw1SKNropcZgZ3M5IBaQtX3MwoXezAitwm88uF9
++lGfWoBMDKFHws6AKom3V8v2JVaI5mLZzBUKgWufOOdpAwShByC+JdNbRILKN6ZiF0kKZ5DrQmC
7JnP/nthhASDOpSrpGeM9jj1nSM0x53BbsYdC0XbQiJuu/fma6PJIncn37e4t9xw1kx9UHdx1Pju
GXF1Eq73QdcIcJm18zym5OaXX78Soj311wTP7TRlXTSQKA45Ph/suGor7GGNbHw+nzxDZxRZhLCi
ShS79dOD4lXcJ3Uoyw6wuwjzDI/6kAPB3rjHTCWqOwh5jwHdGNFX0XDsRO6Qr9MXpLfpenby6MUz
V7Xd3YiYNM9qPYGKWncpcWflqwhxvVfkZSBKs3AUQjfgy1PFvWK5OAvNBe/fYLPwt8jg2ijraGmM
gLoteMPtg4lrc0RPynD53jVLe5w6GZd+ORDsii5IU7QQ9s+DGUUuU6MdqsROi8refF+9GV9tK571
Tf+MmqttQCAmVN466FvRMeOKjzPeSgYenbDdC2uoU0coh+CLJAlx24G79UCqaeUygYX8mCoLJXe7
Npn3OnPLYmUGXs3U9VwTfjREFVnLdxziBj2NNg/F0l5hiouGjggD9/tfZYI72pm5gMkfjVxPiw5P
zsFYcgtYsIRfbfyMg4cCBPhm8W13phTeUvttOneK5/UGj1KrRapc/sSigqA4qhpYA/fzgLdLTPiK
azZUDbdD/keXLkxJN4FAIjxxrNmm79O66pRCwjSBgisBuAO38Y7uJ/TAxAjm6+JTcLnzGLTWMKvS
de0OLKKWfhsTrNNya6i3kepdP7GniNLRNjbs3G8kAZprMGMNj1NzEPtnr0MXi50lFhwFAFYGNmEE
0i1VGMv7pQlzDXtTx9EtJcegAJH6vo74ZjSyfTmxKA+kaV86b4EtOIqhlEb8XKhLFlanoMxcYoJi
AlByOM7/+eDJlcr9Wvo844k9kYeTBUBqU6WehmmfuBu3KUPtBwf3ChjLIBez3KOZgHbWb7i5WXV2
FePHQZGKrW5Lbwv3jls1leqUuux8lKml7klCSyJkzkMVGEOEnZ3JsF9Zu4HqXQSBeYa7SQb+OPgE
wp6dJndJ9jLL7K8VY+DZDtbyKIE7GtjPIGMZJ4MMpSNlicn2sWqj0cxDo479KN+ZsfDt5zSZCuqy
jOb26wJJv3vMIfODvYEZNDxujSl5XViIaWLZ3k8wUZRti88gy7KqQJDj460plCFbu+mMbpL4C6d3
H79EZ7p5tsnSObiQQP6XdQGXEDKudo0px98rrRcFsEuHkOiibl3Mx3sp3pw2QQ21+9Ex54X1sPg0
GAx3QkiJ6nYQnXm1jpHtC3Qnr0DNrve35kNq0gA9+TBS3H+bLIqV3d5FsPXWvEuxFLuYiO0EYwCV
dEmzNCoh9t+nOpyp2n9FI+n4P7B+rfSdbZc4uamhDHK5iHyLtkoiyWJMbEn04sCDY8o3xJmUnOv+
q7oOl3vwmOnKEI+zNO3Bmmmh+cGpQquzUMO8X50tSfPVzYDHVAQMaa8FuNjaOh16JaUEnqtuNcTf
R+HhbeadS7cB2TFxG3dRC2yDxV6jOGN+a//SgkMRMLRtUf7Af+VR1wqZjDWaGF82crB995g7UoQD
v9MU9LZB6YvEpreLUCDkf5FDf/yIUmgk88gM9M1YvQbSCtZ4tcmRtxPdTu87SVKgd6o3rf8Txn+e
RKTa0oSIrZn5YSOAvVvaz4y32lA2V4rrS7sv7YURYCuXTIwLd9fsdCEFtofP2Tt9O7APCfH46C7B
5/P7ks9HzYaGMPkezb3XrztwbFrK9uwyufZAMS5witB6pBZ7D0BX3QA59UeZ3y9MQ/zRipUbhXeY
gFUA/sPSgbVoBt1apGgYmPmmNYDPoi4EFPE05+PsrGAoWg8JNm29poYMjso9hGEjCQcMQBHXkDru
5I2qXJpgBFReVqsCaa2ZW6CSeuJVRf8kvTmyw3WpmrL410FL4t+9g0tj2Gyf3DWzHbgstbv6bb6B
rwwRxX/pWvcdDTMXjxOaPBfwjDYlphAr1WcKKGpkxt96lW+feknrWJ9thr21eFd8pIM8lSLTt9wz
YzKStN2BaNIK0kkjsnPcNl1gTGtPuK93a0PXoOAnp4bWTADJjfeDMS6Kj9zkDWiMG1rX7kWX6hOM
TfYEfUumeDIAjCJBQs5WQnU4oDfb3ud6FnsSItIa44M1MUqLoTR7wcwDHS/rnObYKT1ucg+berR7
r9zXSOzdVAYfFxhnShRuj1eVHBrpWtRoeDws1CSZrqQE82YBBTElxs7wlsgMgn5lDkZbvEimAFGy
Md/uebI5gxuPvJbK/zR3CQDeRhdZ/lT0u7Hs1ZEKNqg8x2g6RpPO1Chb5t9Io4jGoq6EnnVl8VmH
rtcqnx08rvHpwNWKwq12d05BAnEaNl+KGJqURCP78KuBnKdfKQ9f6rd44Bxc+Fy6zpgOjNRlTdZj
3iSg9DbQHMbVqtVA51ao19O8T3/3+IUhZEIIygaLNchtcc2OtZIzC83AyuUWask4GSvSwKt93t3h
YWgTyUsc9DH2wnqNBxhz5rYAcaPXADXW+BY7A7/WDmtobMEiKbqxWCAEPAnlo6klmx0h10gsYuxj
sVbHBJ8Xr8qmHRLPci5ULHEZmr0pYeFGf3bvmUmTFX1XmRrgdc8iDv4anuCMSzV5AJs8m3Fo+CrD
Zjeoue5xl+xm8K9E1/EuhBsLDWhFtqty7LUJHX4zyNDrSJ/v+O//mpRnZtllgHQNHDH4z/aaeeOg
t6sYhQ42mNVeoL0/yd+NwATF282kKPuOKlXuaArHkWniOZQQpGIs6c+FoMgOr+VC2QG+h46YKcxY
v2pkwHuFBoF3pg9CD8enpc3OCPFMzh4BfJ8OEpGHGpGXxZpVwrlGWCb4MweeLzBgiiKna/7raDz4
kuFK03aT0tO/uk4mzMwenTo8rqKyyPfMpHTIOpzURoO4frFkdJpx4z3BGf16ChK7W8RmEbzGAZJ/
cntok2sETG6qHyVE+m/iIsiJ9K8uxXsVCBpwA5joTItpQokgp8idd16eClAMsQIbdnr21N397fZd
3cGRjBEk9lH7L6HRbGg6lmQzA64tBeQskQIWa6iLtaRRNvCvQrxrqiSuDepljZdPWlzh6hGvI995
iwzeBskrtUnxMqcIWT4EXGrqpk2ICYftlAW0RPPm7Oo4MIG83OP322AgwapdVQU3IrA+49S1A/lr
+wINlO5jxhWhLMYUotSwYFGx8h8MFeoqFafyRc5PXv0omfxsAUnYUJciT7dDMZ8Mfx2/rXe0vOv1
8eXfCf6v9ReA3J6GufcEf6Kgy2Tg4JPVEivz4OMXjxkt90wPiksnfi0dWMcAXORb0FLirZqDOOuo
uIdSeaq3Dc1uOKknqMM2m5YyZ2G4u0aurxa9O1WG979sokAfM00riuX3tvWg4+rAxECaY/mwwVn3
ZhF8+vFMvcnn3Qqn0U+ehNtX9mXKrGFmW6O7NMqPxhRLf2OTN4EEX9lPFhoVpItUUIh+Hai3ydGt
82PCVkurNb18rFSRHdioZ8HpvfGcNbjIxUVVPm+CA42w4QiZ6j6xrNOApLXilUH6Ena/sp3vZDP3
9N9VYtYkwfh391pUNctXDUvxPvEqjr8w1t6d3CVFDBImOr6BHhCMX3NO+Y8UE21tm6XazE0KDcD5
XIRfzFJFpwWpk7Bs/telWaC40pf75tM+PcZQf2VxQY1E5dCOHN9iPmXGYyafboHbZMRWljMi+VlX
Km4TFZAWwnJkPUczrGO2bvInrvf62GXPlWYegz/f90lnO8Swzu+fOucDojpiFW0bBO0Ynv2QMOst
rJtCA+2qeUKYKkjMExjvNjgu1QZeWAPfxOOkLlU7F632sUTbq+gWopxDKqGMxXnJvD0u3Pp/wcBI
r26qSlnI37iaKZX+sDnjn4pdyxgeax9bmowX5Q7XiYd1i0ONZEisVJ4O7eBr9EXPqr0uAsoCxTVl
EzUWVEkRtomfTmUB9zR9dhDCK3CtZ6Wb+yjwmhIQu54An6iX/1pqYLpg/qqJ6WA0yWeLWWKoqOgy
eQ32RkX7z3L9ghrI2eNGvcrkOSpRgZFCxWXEApRJUYcjCYEd1pJXlh4N0V6oye7EoD5wfOYKeovk
y5Z2ml5+KKGgGpGWCUVYKyTZvlXTMWRPkIef0a7tu5Yp7rFCukK9T3nlXcIGFUtM+3wX4Xsom4fl
ujkSi9urpMgfz4gpLDAdRdBVLuX77d2RT0pOC77yaw5Atth2GnjcMtVA0Bvkq6dwx/FNLziOhuNv
nkG0aG9wq6dVavor76ces8gPmdZ9c2Rq/IMqbvaH4hCJqMKKuUIJVoj3USrqRt4Xz9CocsZOCFiN
+GGhWrHALLZ9y+MO1DD1r7+R9VMnGnmOR7xHucK+sGm+M3QlXbrZt+jsBDNemcrxCCjlTbodTsER
hEw97zmfr00WKny/cmdKlWnUpc1QPvOdGmmpHOmgnPyibEkYi6NxDIc6T16FMVLh3kaKMK6xPy50
F9kgA0CQwjJr2Fpc2xrsHreJWKZUaizQbOWtso47a2oSUoVdX2hRT13upPHqOQ/BsoRo4Khjp9jr
LNvXlIEDA65iMysldwCvJuzAsv1MOnNMp4+aQTSKTyRlLhr4NYbtcncTTr4pR+j6cITCK+tktda6
SJqiRWYgSaJwqy5KyDeiRTTKqzHrqsX7xk5LLYtTC9OdN9Gk5gs9Cx0jAK4JmiUAc3VLZ2wiYV43
VBmPrrtxGHbBFFJjwn+JnU5YW6hIiIzaJVSHKwxBGUI7cwp4caO8oiz1w8kw7OQGUa8iLp0uwR9w
5CdFh7NsY0pcs6A5y3kJHeiJ1iQnP4QhfOO0a6J46InnuWCKGdKLt/K/SLeMayysEhzZc3y3Rm9q
X84dlEpCWg0gdP3WXQH8hwo0jptZr7PkEnEG4KwZ6GEnwGoy5XWzbl/oEzSxLUJcx51Yp21Tf2CX
FMrxtui5PUp/yN/30PbLBy5DAAnriCM6Qe0mmLcSNnvFmR9EaDk8Po/92AEqOy4er64at6LmlOee
c14Y1lq4ZtoDHSzcdnkAdRpFId03oe3QgzSxzgKQTLDoMvzAJ3vXgUKlfQ1K3CIRJWV+HV+bC826
amXaJmJWv9TUs3mZbFACoYIMUO55oH3L6atc8+j8HDS38knYnyRjAgDFMqwvQgsEj/SDBpLsYRVB
5GZ4xzpXBeDYbA+INAb1sT6dkP9Ud+Cfnw9faBAyLs5R0HLBGVDd7+/mJ/veqTUYicZM44k7eFGw
4y17S1aCkg0+e6U9LygLN+FrsXYeHNcpAOBQUyDaZPSidATGwCcntDqdb18whRWVZ83CxFj03Yvd
ApFtTX299KmELXGZjKPL/BFIabQctZcks3zgYKsEbFQpUNXPQdGGQogKt4GtxTK4pynW5+YH8FNu
Ys9EL5KDQJf15ZAZ3Cm6SFWGK6E4/Ts1cNhNHLnWdBvZMpvNKS3WoXspkuv7/1IXCjVIZ4Vr0Jqs
SHgiPs4+bdR/V1wyVs72Vt/qNNHdAwDEfuSgMhXfmm800TVu3gP/UKvwN5NLfVvxXp+UHMavTn8F
BQwdk606g1uGUuGovVQAqheMDazvA4Y+QIC4hdyu26tKzo8+RBZVqPFQdYRHGbfzZxoBDZbrZjlL
GzAeQ3IKnFe0Jo1MUJUMRRlEGrDJ3376q/+KdeD4kHWdmDGvNWl9CSQ6cq1pzTkJrUAuiUubVbl8
kyIf6LrgbCTl7nXvzh8djSXhC7yKEsy98CUhbwQv29sVMtWkIIGQ+wqtk/WEhvoIcnuct3MfjKaQ
BOBMBWiDzh7ole6kjGG+bmBF1uImKylR9x9R241btoUkjcDL5RdHpWy7z7/OitZL+Os2sPUhrRPR
+JGwEzZa6IP5FZnjHMzMbyuU02dPG1Wx1MMYe7kOuSQ20PVjrsfICb88REcAGfwPxfaIqXNZzmgh
UCcR1ZLsILoQ1wJYFls92hOwlQuv45iwg37+WA7l3XTVPlJcNCHe1L0BLC+xZJwTL9iduo7leT7V
4grkQuPQjReKspyVPuqBdppU0sGAQnL8mm4lnu5OduBkQ9OkL1HQs1ZeYtrcmL4EbSDVfxS48QU3
oT7aHqgybOqt0bUc9rEIHSqoG6gHbQcW0ibV9Jw6IsxTZ6FVefTwIL6PXadvOZ4adlMlObqtqhtj
wuMlGY2R3Dcgwrgi5Jv7zpW3kbh2vof2dnhdWnKRvP9rZFUdMcdmJBypWQSI+/KrxnqATwKx3R4p
eKzwmWQuuDknmzD6kSKrCiFNBXHQW1XASaaUWKtf94K37kgtwIVZ2bfx87jzRBH4O1TvIaeln3+M
9JZjkiqIBl1NXh1hiBPEAFSHt0WjlCA+AVjUgaTOJ16vv82gWanAzE1mh6bqZouGQ4b7+LBhOsHp
G96sPwk/ML67ARmmMFg4edJ2GrG7ovYQlT0TwWQ2YJn9w10UV8fECTa8bwgqIKV/SONoFXlLlB9C
TK2MhgHG5lQolwdxID2i1Mgex2juCcu6dyxjo7wkZ1ZWsdfkl/wFquuKj0G9fR0f8Zx94ro54bBy
KN/ptCCmrcJk6zyMUAk6uofrHLn9MstExNJWUs6l8/Eo8I67F0VsLT8ERUVRHY9ZHI1sU105fYbD
SpphKVTD7RGyHLDYL1GcSMSB7xCOkCQe+MoU8pJby81WocwR+WQZLOv1Y6PgnwH52eDzYMG1wMJG
QHdo8Hd9vZ6yBgvmPhw/1/qaWkt351HKnX88YxKHMzia6MomgA/2fIyeaeXTyzpJpjCM8NnZkYKw
R4nj0NG+IvpCTZWfNFvEv9rI9lRmjEIlYteuHm9ct6zYRzclTSNK7ggnF9wPyNcoPdhuP4H8clDY
CHuvyqnmNPzkZspS52tBVY00RJTzzf1MjIkoD9R0VDqNttoMZ5P8/b84LHBvzz0bXIgAB9x/2FUU
vSDnzVD14eZ/62G/54cyYoF5+tiCZH53tUaNuFtly/A42XwmsKURUzvqkLkJH7tpUgPsq/lA4oN3
c5HE7eczcDu8TsofgLNJHuqmQ08cjGlUdlISXuEhLDhKsOgSFsPeQVNqMTsdL/pv1b7tK96k3ACE
9XaicR80VsmTIN1XLAw5Sm/ptxkxHVxp8cw73zK0eeXznBtT2wqa+3aIv0khFJu0jB+YITMgpWcD
lHRax8gFnwJ1lczbKjJEi9+kXn65Frt6wNwErpc8BLJzl3ArJJklF76ZRfVeROfHEXUYwjz/eH9U
vO3hg+ez1YQ8AzZjlpf0awxE7Wt1EP8EnAmL/gnWq3sWz7chLVhCf0tsOQi+404QtcgSagmxiqzP
9TCFTBgh4xyfkJJS1h/eb3SHi9P7hfT+mfIAISmEUNppM0KiY6uH6gepuanwtk5vp9Zr5az/6BZm
/WfvYV2ZSDlCTYLAbjFbyvjs6vTw5jLP1P1dvbhV4CttIKHw8NlU8lmsTNvWaE7zi/MyBeKMGIEr
B4vufSYLDYyEN5ZOwFzVgSRbRoKVGt6ywaSCLG/ya6yocdyRZxG+7TK/Cq7Un19R7/8hIs5njcEt
gpRgO1X1JuJZn5BO0m4QlM9x8hJM8jDEiF97PvXkz9ckhhAwvhDRGT+wtnecFnVODxWmCnUw+A+O
bFkccznOAj1ox5QiSc9CxcsewLX5oOwscZJhyRK6YZxGrX7Nglps9ayIHyNAkdObqrA7MLBxC3r2
SqToksz16TUB56i9eatKihsFWsh0TuXsE3yFg1lqp+ETBfWix3hPfcTZZjJXTdrLu6wi7YZndIJk
NVDeB2jKXgWvqej3qT/OIkGe+V9FYRV3fcmryi50ByP9HUU6VgWXYgCpQhWDz2ron6stEN6EtG4t
zqe97lyl8evlhY9FwUJcGGkUo9LYI0MVfKOx1hxSczxgnkBUtqBjtAZmBynJ0Vcxxj/aaCpHXv1I
tAA/KaHPLmeNHDuMTQJE/hNbnFYwSgbuPeF/Y9OulL936c+lQWX45GgY2v4SxRDl2yC/eeB0+eX2
NQhKWHeSRwdXR8WzWf8y4pW2XHoz9vMvU9M3PAICGlcaNPQud61b2jT54koZ5Dx9krVnI0dZXyYe
Z/ClXEhSLqKpLrXgoU4P/hZE6/nRTAYpplM5v4xnD+Re/b0ez+q2KyTMBswMxW6E9kHCi7jdqHIP
yT0Ruqv/in+OFCA49OcZ0KPp3Pupzxuw1yoABOc2E6DrgNuffhkwQCiOkk/IBHXrCYu5m2rt6k6G
lryktvnGMvtlNCkf4zvJ7TdPYDNl9Yg6aDS2n9gWJBNZA/zFdq0aZNgyOoLzn2abmPqqktxv8K1R
2aKhXOPsAMseQVgv1j2gdm65E++Uu0CHKFC9Nudzfcfqu3TVH5gn6lCzGc0bj8fhK7aNrE6d/xPu
Oa8Vg3QYRGO81D+v3CrJ0iXsO0wp489AkMzLz+HA6YAMnveRJlhWh0awJS955nPVGt6NS4NYZ8hw
py/z/imhDqJzfLrL3XlUlr+TOUAOoGTfzQ8agERo6AYwj4fSNdYnFxVXy41lu+PlsiHzuVTcC4Qk
EG3efFL5DWDwo3e6M4BHuS6WEky9R1PUUWj8CO+2TFnD8Y6nSbOo5tjDXP6h4Bx7c4PSfKiabaC0
sXydQ8/0hDpKyhE5ILLa2if40E8GDiyYRGfyZLHamUTPp4g8rFo8SNlAroe7+sXV/oEROHB8cE1Z
y3fHgBXJvtABNdqwi3fAHdl+zDXARxjMdeFeRGMsldrA8oXprPpcUv7io0uj7r5exoJA54tu+xc/
cikG1200GawrdvuvULiN9R6TKbhu4GmkTarGM9qv+X0P3FU8jTPs3UFK9hIgoOOYYQ9vkd11SHxR
Wf4BnN86prH2nZzVosCqsDIsYgJG3gWpVrYA4mJY5DW1pM//AA+IMR9pMxzBaH+v4jnZLxeNfPh2
9I8D5W8WaHpM94D2qjQPY2qECd3vQ1qWTMR03Y2xBRsdJuHA+IO4SujDVIFmkYsfjz44uXHXVMI4
ffj/VDjgByvtt2FV+KQ0Cu0quheVOFmKR0LW2rBZSl+0pQXegqikXZZYfZFnno/FwnWtfBxaRJIs
UxPYE7yI4wjeTT3Qn8Y6D5urS+h6hKtnCrkzLmj1knF4jYBeHJ+kE2eyqkyo0f4YICvcIv443+Lg
IvwUPZ64DbPBbhh81dYrft8tDRP+vD/MXZslRmizd5CAxRodZLOrmJfdB5P5ftziaTyaUCuV1Kvb
8RnoFbW+WCSTomkiq8QZFzoF72QWTIXS5sj/m+M/icTfVemGYDzDq32so5Dc9M9M6Lc5GOh1t3Uf
t4tbgyvMtFWT/9JriOFq+Fy36BkKX4Ru2K95xCuyO11qNsdMWjhaq3KSyf7KX22QPSumX7+AW1ta
LF02eCTVKZWyMyrLgNzfWjNVww7R/qrFqh/b/gQXsTXrOJblvZA6P0hCP3r2JYAzZ65s+pX9mMHY
A8+KG+td35g9V1GZrDH/2MkwBXeGYW0FLRySdxeoswSbgpNZslyg0UdOomz1zCtghknCY2KbNOtb
AQpQmy0tcqMZgXMJA0Fr/WeM3c1ulXZY+U6tszEC5x5LcBjWaLlzPGgav8Z0tYLnZjSvEqJyTPM0
7RPaUGBBYuUkpqTNx064Iklnd76xea+FAxYHAy969an+zmQ9lCxaQPYkWc1qkhjHf9CcTRL8+4aR
E4bq5U4UInarg/u18xTg1XFhXnSrzSBBntBZAj1Y6AAVePt48VNjQCqfjURcOeJFSYsRF1i8HKur
nGby0tgdQSanKv5VMQ9P466A08qQjEPvtx//bhKQe7dTEUrwakKl9qq49dlPWid3sVqPvYVikBwD
BOmypj/o291TScHS9EJrwKHb9QtOU0/0uH8Xucyj+Yhd1tVOBl/3qJ9G9BhMizIPZ1Zv6iQJKQAd
LNMIFYvDs38kld8EexaJehB90h8KzF4aD0BYPS/l8e1fd8b8/yr6vdm0ywPZF34m0yvLxbx50zz7
4vjvxW0q7aOkJg0+OZuJSv8OQXYUsFOAqaRwxuTPWyLyh9/NwlzSp46m5hFWiu1Hj5HAof1u1QPv
/w5JFIJq2UtYvuUBtiAaiEVTcB8clDV3xoLoberdgE74Otdd9+I04yHNrabgx2vBqc1Ya0g/GZUH
xAFtV+6+wvSM8/6Sh1dSog9i1lW7BtnKrXzE4CziBCAaAu+6hWHvwE7lAZhB01J0hIV6UXsmihqH
WLF1oAf/UrCzEycLPJJyr7EbEu65N2xgCHbhAGP8xuLnrDAv/76kWl3cvTKFyKSDvKy92V6haLF0
PUaiLScQe7jIM37UmimJfJO6R/Hs+7sbeO/dgxzKICd5P8+ZMqkJXZd9vboVDRUnZyeabcKDpoVe
D5WCX6nfXsQzqpFVyYYMGbpZ5/JO7h6ln4wzXOZ3fOCjGMW8lKYRNEnV9zJikETw1WgF5fdOVYrn
haW/2H+KdhSfdPzMCfndpZqKPYsc9hJwW+5r55ldkFwknMkWbfzYD3dzre93E5uhsCegqwVil9Vp
1vI51HdqfmQs1p9PsioCbgiJM696avP+AlgVt4mQzl7SgMKAOcnZBQt/nJYyhiTM74jD2mtmQhux
yq81rEEKBuZle+b9dOTmkGPPBO7Ex2083HzwUEMS4gBOo7GF1mMYgyEVdHByijeDHvM4amErssjt
TEBdu3cUuihqN3pUD3HxBU7BPoyHeSb1XgzPSPjIXyJGp4akLd8a57XvKNdAGCUoDj7TArrWjzw1
wkcBvH145BO0ugKE0GD0re836iAMmi/Aj3yXv1TUmAJevSrMmmpDVQnQ55Milit5UEx17/KJFPbu
Nv+lDec7/r2kuk87kjBP9ZiXYNiJ05sKyuDE1QgHl6h6HTje4KhQpMdx/R2G83wVMJ3QIaxR0ALL
8ysNcBMztu5+0vjlS+/la+EQ2+3O22Wg+c3sGL956HR32nUP0NVpjbCou8K1H8DCZwJWukQ/maDe
bvPoO2RPAkWzA+KEV8XY8smpslL1Anmz1Nvo7gBBz4jmv4FuR2UZtyZUbt1QRs+So7PWlBasAXxL
SA+UPHpZjm/dHKGf9z5DCC8TLTZfTmXzCsiQPxQ+p/GF0y06cLve83bP2phfCoufISmM50MTVAMc
gZppDYK8cLe+ZQJk3rT3VuhHeX4wPSqZ+ov0LV/+Zs5fawGU9kB16aKXI+N2GSnfIbpj0Egn+7ci
myricyp0OijhzeVzQYsXS8p5r/XgOr3OGUjxjTBBosgblHTGyBNs1O3kWHUEa/W2lXlzwI/NDRlz
ISC1u7x0dQTc+qtzCMjSqpWpj4EcaTTndTJngEP6ew/2bv4m3Ppf4z9xFC5db2OeAZ1FgplPkzr0
fpavR08Bzz16hxL+GCpbbA7RmepwTX7Lf51L8yu3FlKEGPiZFXgVTBtIxSBnE2W7mCVsSnkLF+0x
YkaWNjUmoutU3/XwGHuPzvgy9RE9VvYze+UEiAOloAx9EYf+h4muM3Pg3ETmghiDj/qgxdvQdpG6
15ZaCxy4+LO3ObukhNa9B2cCohs2ounOv6kWzvRBwN0JCySRMaxoPtqvKWI80/bGqoYvAaTK3/Us
XHpGRkniJwG1GRL9Vs7ymKLLFBTqYf5agAECln8PNwkwe7g3IgIbGnaQu4zlaohOy3nipvASQAhy
2EBX7Ox4K5Y2Dq4gzQ/9q4IV2rhTDJ20XUXFXhCkFVLIfz74ukNL0jPuXB5TKCvXosB+o65rIFgi
UDrSdNvKmrERvsZJsDYkFrlq8rbXwQo+qzwrzxvuB3wzTJXpD0ztAzXmXsgCE3OnM/9JCvfAd5OZ
TsInf7r63d2bAedJopvX/Phw9an8rtCyVA5WAHy7IT/y5akQmaQP/wWHWX4IJxWj0/dHKTJ4PoU8
D2FRoyG9Tw3KXTHPgCHvi0XNV5duFbD1nag9oT1pKhh2LDDIGPfn8mc+YntEOAlp/t+x0xZoRgEs
TmupWwFUtzUALSMBXCIrG9KDLAvivJ+pOO/NwsOTFoqnJyn1hAM+HK80VUtIJkx8H5Z6XiJsHoEa
0m/k1XwQF2wUVbHkfzLTL+tEyxFA3a9EUd9lXTgSpDUJZJKiVW4Yk7/vbEHe9O1tdRsBCr4+p5o6
xHtFcrfJGd9k4BTdaORvBqGu6q9jAsgszO3F+88/mEs9ejZdZ3FavXPpa7fj3H0rkeSgbvYTUYcb
l8Rj9YY/NtTD5ZwDsAH8HbtCnPBMPQeRMnSkD1hpbp8WyZT/1Kw+TC7A+eyhXTvrW57qz6VMqLa6
WBAs5uhcsyxrVnVnFU2iOOoDDk1zH6wGeEZ+0w44MdOnEGnjABDoYhCSdRikxXOkkWtQEsfokCdk
3xQadm3EwWK07aJECX5+2lU/o/SwOoVydnwLoqY9qvWHh9p1k8+dvVNZIBzq6Uu4L9Z8Y56cL1HL
wTCyRueCFdI9WCST9D1UdN2aeLE2P3OljACt+P1T2Aa6OSgLJuE3kWPKpebzBI+2ZhbmkVHLA26R
WmcUDPAOxqygj5hhKIci+vX8TJZqPWOiGknxdkn7RpqBeqR4+Gijybl7L2YKJ30nZGS9OG26eX5E
EcL+av8XBDSTxTxkGgo5KUDxFIQzo9IFHPp6rpaOOHP60NyD1Wcq66dNMYRU3rTsbfAOdvvkhEzs
nqAplFVYmn+c6MydPn3dGwKXj5gbBL58NRXdagGsH6zKaEXne9CTI+jYgDAHl/3maNyPnZPin0Fd
llv2xFwlOcnPtLZFALLcZ/v5/lwPIi4wUtOqqJTw5ZLM6c5dAENiX5eXnyqkGNxZ0dgHJbZVHG/M
2cnfLkLCbcYojdturFFokkOW3DgWovj8aSoDeIwZCk3K1irkdVf31HXFTzzcIMAhdcYlIIhfLa90
hz1Dgy34EtHQtrVGN8qJmIcuvn1uCwwvTq6oNFuDYjc4gB+Y9ivQo4MLVTIrjPZQMhTbNXsiMrLY
LsSVcYD7EgaBIOAU6bX5NlpMCeNV//vJvYbw8JbGtORj6UGS22JGXuLROvJOMIeiMs8mrogLkOk6
npzsCDmBTP8hMU4FvYdnw/r+noXGze2QczCc7Nbx9+t0D5c3hr6OAfnky2IqFGvHesub7/dTCDvo
RI7L+NbbxE2WmkAYJ29naMKAMVhvoGZ6CBLkucEfbIP4bktdij70hrudUeFGr60StY5filUCswgE
BR8RmaXibGEcnkx2XfKyTUHMW4OOwF4vJx6Mj38oEk507asdo48ZFBIGSBkhqUyVUisZWUmCzIXy
WnN6xaLS7aBeDz86m8s1fJgMvDOONrdLz4m2intZC+gyiAQyFf2HQLzTYpNgwryNwL7Z9J1nvJIr
JKgEHAA+i6nc1UD/FtgGYz3CLxFadrYRAEh1S4CG2EiheTzLYhVsXxjfMslKP0zWn1YAkux+cv0+
J1+/YMDCjY98mNnvk5IMGPGXJHVIVS+FkDTNtkq/4eMqPoym+9gFSmWrNETEi+/xXrGMdD1xhxIm
9TtsgPAFKYiBeNZ6aDn5TeMQDxyo+EW/VOBZjC8uYCNAnYUOXzYa/jUSUWFgRPgcpo1h8AEzMNSa
F9ktwoNUeM5/tIVzJyFfxBaeQzS5m5KwgG6/lGXoyJx0VWlafqzIOGeUTpQKXs6DCSeIE1bI3bTk
S25Xeaq2GNM7fFO3t3bFgBwG9yh/PD5ZMe1PytTA0SeMG7S9wdE7XqMD7Xu+2qTXiLAl6QRzC18S
S3P7BQx1Ng8TTgBc+SqRRFdEKczh03nrr8z5cBYoJg6cohDJws3MTCrFRfh3X9CuNClPH5XTnrpP
Wah/4tZXt70V5dp3NzMH1r6/luLVzmecESK3TmvOOlMS3zP6uGxG6K2uaNW8ikszm+iDM2NfH6pn
hqjfk5hOK29CeZ1XUY+vC5p8/VCWLXWrP5cCyckE+wEDiq+DZjMUMIKet9y3WP2ykaSuoJmT19u/
b22kCUcKU7FCDDWURiFTUgyDl3n7o6YJa4gDrgp90TR3GF67lRoRB5IcFazruMEs7uzq8z98p4vO
FQBIORzdkbi7o+Ku4EFp9EW//MuAzWXH+kK33b30J5J+i0TUQotpycUYPPnlOCR6R/TjWmBw630+
rLaCZWZGIFmU1h2aWvVCWKkvN1oZsgQZnMh9EvyceAFB/HBoQJafC9ZWt1Hi1p7GZa1x69BShDj+
onGIAMjBNOxsNmcNya+gyAP/6OKIxK1DW8GkvsrtjPcNj9qLdzgx6TMJozzVwD1O+ts/TjWXQAfF
F1CpoUueiej8IO2SEdBeqGQgyDmuMxOuwJTJmP1uWPF48iUU4+q1kfHGbVY8mocQbProojVw4G4W
LCfkcohJKBc+L8T1S2jszOht2qxi/De5tt+f+rTY5WNurVNt1aenTsXuiMtnCU0ZkZNNFPZbh13C
DXthz5taxLEELB02OwSkzwtMzGYsbhbrABGSQM6aT93Iv8Qou6qFyyF5NNn6CycQkjsUPwRso9Vn
xhb0gdVPQy+f9S64TGcedegLjDTegoffYwBf6o3FiIyM5usgWKeFZNOVKtzQge5698gyTVPePa57
5x+6tO+QhBk20a0b5uFYkgiLKD88O9pA/F9hNHia2H5TZ7+N+dMryo2BtnxrHps3+4YseZPtn0n0
zJid7jotMLSMdJeUZTspdwxfJsJcZZfbLY/b9xOLcCxjT4Qmj9WELieswORN+qoL9SwcXxUgSaWc
J8JI0J8KV8w3kfyBV59qHA7ES1jeQifCUtdc5YFhoZFWLSkbmxudeX4GAKunaHNrciHh6j1qEOyp
onr+FcSNt9Ajv8A8Poq3PE51d/sPtG3qSRWxw61uPORGRGpGfTO+X+7mNEhMtIfZ8pWbrWUVebjK
gEnjrz5AvqBmROjEy85h0v72Iqx+EuF6dBqA4dR8zfG2mhrNUBg6Kt3bvL06np6Gvx5zuIEqCrQF
45wJv2e7O4MEWbsVj3IoIfCi6LqSlkVhbBgx43hI/YHxvka7maEUB02XU8JaLeWGqOfoSjfRMQbu
L2GrKsXO+8vDwJuh0zAYDhXkE8Vbx+DuD6S0F/dQcX7rGgPanRRWwoixEAkJ5VqE8x8Yopjlr6XR
SsiA0Fe9OWuDZCYTpNSBaXporbmTdQCWTLQxpwQvoPuQPaWw/yPCdtN4VgAyStGEJqSwgjzIwcUo
CPLHYv7JjqQWXHmd4YD0pjV7UUP7tWfZQdWFbhShot1NuoX6XcTQUjokz2oh+hzGqf/3o0APslbl
ZusgpWd7RT87i27IayURowIAU++oV5jGqaG3iZQ2YOxbIO0RXmXzXBRyYFzYdXqzL6QAHkflblT6
SAwNZNH8zINvhZpymuQeMrq02dtSqdpECZ6BirED1rrUQ7/ALQwD0heUNYAuz7VEQJy2VdeJyoRW
OWQ55n+IupjU6BgIl6YmBunShtcC4jAqgoNSNi/B5Xk9m/kXCgHoOR2orCiGu8UFQd2ZAnC1a6xt
KDrDhXXHLGP/9C3r0GNB7YCSIt3xEmXvOlS2a0mR7S94/oNZditK6nD99mvHMBgAGYBKaymkqUDf
+wojmj69FZtbaH9r/I8GE87j5DkN79Q745bd4P70+nsv/oqU3P/ut+/Jobw1W3B5f6XOvIlAc6Y4
HmmZT6gU5B1768kEFdcRTiNnkmPktRNNA1ts6MeHKO5oqYnqJZlwp2OmYx8YMWakaAHhG6A8qMra
dBprIxj1fyVnLPc8JMiULDu4QQLWEJZiBksd0WBhG0fI8j1G0w2GMVfFP1NLAa0ZXS3ztZZCKc4g
qtW9psxF3ADnXY+TlQH4GEwhKhODOd3cb4GpRR3wk4ntG4ZanqgrtBcJ9a4BQDX5RQdEt19KR1nc
YXdOT6mV8+oBk9lBA5Vle7q3dvkCbXN9N3O6ItTLnsfEhBTEwnFP6k3YsBy03LjTfqzG8db0pXJZ
zB3L4X9sB90bzYG/pDv2oCPfaeTwVVHEdFxDinaZ1weAgA2FjxiG1NUaAsjrDE81PYu3tB0ZoHHR
y5X2AI6BVzd/OUNYVUErk/AzbMRAX78AI9Hm3pR9sZ4xsyP7UtvgAvDkSPoMDYfkl+BtbHku+sCw
q4x9XHLrE2fBmgypr0XDdk858Jr5HgkdyP8SIQoPUUaYeUlnI25k1le+M2cOvOT5Uhh2MnieCRtG
kmf7cmCCuFOu+/r1YNVlY9rTAJgBn6i7z7HluQ3bab0++ZrXUZrg5QLtA4RzifUbQF7OfKyUXBz2
zPbv6TQHT0w7bnP0R0y7LNQu2e/0ccAzAXaqn0jBfsNS5vdDkhOMksrCSRaLb8SuE9V2O/1nqlC/
xgrV0zniP89Rrjkq67oI/Iez4VkgttWi+ZGq20olRcvk/bnJ5E2kqXFUWkS/InycMAewySpkaIoV
KJq6R7uGttIkCktQCDkyy6FXnxtQzwA//3uA4USWPYuKcDgg8kOpCBSoQO9ssp0vRaELyFpXik52
Q3XxTHsaDr8Ik1CQQatn2BsjNAqriBpnh2heeUVjdPg15cvyIFLBXdUxGiIF9spdbjYCqihR/98O
vtqinplU8JRmz+BRSQDg7ZzyDGh7SKNUIUjsGjy5G0QMs6BDCbEv0S8WPdXR7wxpnuvXOPU+FYfL
kvUIZr6gpvlfmumtUzTXGOBRH5WZBUvd/cfeLoAHpuNQ0ucTzk9rXjJabfAUEwck96VC/LPbZHLb
v0+Plo6ciVHmsIe/LyQupNUQxZrie3pJhXxvlM052nJ14feIs65pKu74nxPhlRYSK698BYnPrYB7
sZwJA1ERSdSwR+HyHWZVUe/+XKDux35umaaTzfuazV2ydMHNGR8gc82EHLACdGcnWXg+GQZTG5Jh
Gc5neF04kiMnmqPW+Oo4kpDWijCDhCwkJ0cv0888d/c6TWZ11aet+kOzVtOu68NGvmPrDhLAtSsd
VJ9BWLloMAZfSoXhJ1t9xvEGT7RMflGRgdPBd4jOrM3Dy0CsttjCxcH/9Rl1DDA/8ic38ZcaSUiY
HOHg31rcYNtmcFmhb2mXQNh3DifCrX6fUuIMdZaX46aCgcDQ9jqdznBRxV20wg2lTolj1CjK7dPA
Pw2uthOmAAgLCv5ZO4bR304ke14MY1o5KNcojwv70uePYoj1Kh36HQfnvcMOtLjxUd7fnehMrECl
5Gq75Et3oQurRxtaojgG/Kipk7G2eD1qOaw85eyqs09a6mGbBGat3DIMv/ZLaghzRxYXmBnLZHie
wKRV0PCnxATHwNIYLHfupWRrbpdnOiAK5G6sZIcHb9632HgrlQraBP7oRHyzGysHs9ytHsKp+Q2L
9Ej716EzT2ulYdMJvQwsSymMlqnFah3mMI5co4y+IEOJrZQ/3Euhspqtdz8RcvrvYZpEBgTEVDkR
IpymGbTc3uyzp1WB0g6DG5F73dP/t6KsSFtUnXOXupoIkoW4ELJoVSIc+O74hyHoPSNLVS7fEKtx
sLYph/QBq03E7xj1RQkd13lbr58FnZtYRuZOhb03jLwxZA+KraeI/t3FBwDa6u114uYOZJ3Y0kPN
XBSuqL8tKsXwrIw3QDg9qhBdQkbg8Ii9scFFXUWVWC+uOCkYxr40DSCavRp3k/7/qR1EoO/Q52j9
u/h7z/6K+GNCJfGLaaJiCWXDIwIIl1J0IrVuL/+bECVckvLM2ytaEUsTP4uZVPSQOW1Mz1omr4YC
8xd0y1yHyLqqyP+JQL91ljWOaobSxLQ0x5RhENN0/FYloJ+EpyFd0JRQUNVm0w/IDfBB3V499NU1
kXCKcyRBzyHV2R8BUu2Ny6ILsJ3zTHZj/bXQKcRbByxAG1obhfpKtAtJumkeg7q3siFJFv5WeNJU
nt7cgpHvB3WYLK6dAXwYswv9OLtO48f8zWojKJPQqw0g7brTiZBXx/VwoC94a+hwsF0S3LwsL69U
CY2dpHEErQ+UTrlD55fpwl0bokaPTUw31EZDMLPocaHuorWiMOsEkG5OgkdsBTjvOdVY+velNv18
1pSZREKm/iNVUrNVE9nOkwfsQRITuBsq1kI3qI/Sgq1RMa7E6G/pwWlZVgKoMTofd99L8jGQDLHh
p1OkktCl9h07jU73Xet5qwOVPJRfww4RpWW5TJP2Yl8vs31xiR7RSZnCOtRJ0EVuDG0E25ybE7Hj
A4ZP/vIbr3iI945ZcvCVHwB16EzuUzXvyjwdNgrQl2oOlIj8NjqMNp4RdbdGjrsxR4FhDejrp2va
7PzYQ7m3eD/7EbcSCSZh8T+ewAjEgDLD0rmLWKFZDW8dwoivoC1upBV3MxSKGhhQ6tJ1lnXOxT78
9TMFCAVCtuuX/TBBcKBlMoAATbQJ/Ke/v8L5i9Hhjt4dj7cxlBSDXpVBwriXRoFDW8tJ5WtsnwIV
jN0V8UtmqWXaTPkrPJiMUcQZjQJbg01zipR+hhYGBIWicE8TfcBAF0dOiLrdn5r1qWIrWD00BTX/
r5GARFZ4OUW4oUsVFjROdSqRLom6OO0gpPlVJqCm31rTrkGsWlpLhtHczI7QxuylYQekBWqn3Hyf
23ce0AV5eXP3m38hF+WUb31/TocWQwLFkp5ktk0rpSjgK9UPJwhKd/2ThPqO4mf3vDsWbupdOxx4
/0GKN/4NrjpBc3bY5f1BTsVKz8qsb90P9wdr9vyWL6SaUwSRBYdc7vj4QzKA8IKi0e6AgNRx7UMD
oHgWcL+4gsrpy/D0oW8jLNG3lNryeVx8GDWxbIpuUO2K+dyXcTsQfRjLxWMqQ296p7x4+IOrsrtD
IqoT1o6K2FlgxC0cel4vm7emljcaGpVwZRsdNRxsGhuqkba3A5BOGwox/tMK20Pfh/ArY0ND8S5g
fjKlWjnlrpooN+Yja9dAvUMIlEKIDH2GiHKyWOhDx45huPORojxEfT3XEW9dsgDSWabi47ERqK0e
WogKM/fq5DTd7FsBD5Svcpq99C3e7s6+CARpEkkQYP29U5ZK6L/ePcwOh7hTe2RStEnZY6i9OSe8
vxFVronmiiXnoK2zPQRZemYyU/Bj591ILAFr1gbqDmBiovNOImmvIx5S72OR0ucJjI5d3lbzJmGh
iPkspaRP9LF7Lcda57M2e0V4cTeL4BN01mtcFQiLU357z8sUVU6rPZxBnIuB5H75mfmYDLvTXuBP
F1koo3FzAaLflEcfIHjbGwuhhlPzoSEPsBJ1mKy8ZHrEhGd+RcKaCP1B+L7CpIMY5LdbjX0ZFI3B
lEMvgi4SoPvRUVBMxT317Ay08rFr+dIBmZ2957o0tCr54Q5odu21WYo4axxfTmg94FlYtUhF4/KS
HfWEAu3pUUpVq6Jcuo248U7dW+1dhOKbjzZjKvkuZ1HxY0+6ft0Dhpzfrodoww4INR9STU943UcD
Shi75BDmz4Ff732uqd5gvfZO/H8g5v7Kd3Ul+fUgLL0NK8gdf+T6tFdVNDqRfUL6eppMkh9tqstl
wXXPDDIbZOBYNFNB5lsgLvcO4uqfqguP1RvzTTU1pHXXYBpFvUbobIp5UvHJzP6YT9MD4p65fmnv
1YgxfKS+ErUDvgZ8gNKJz3CQ1PktV3iwy+kZujjiykLkL/BusweiBFDBVaqmQigGGaf/DoSV41pO
sSchzYzp/d5Z1TF/NoxDR0FNSzTw738aKGDyqX8vLaLwCwGa4uEiDw0LO4T8U3etb8AgA78GQG1C
7C5eY6wVgw6cIwb4E4y5JGZNS0uYx8cwBZwKNE7mg+N8xvSJFLI8iSB2ZWB1ZPJ5Nap0smpLWh8J
u9rXg69KY4meLZj8ZKmlbyu6nYH0Yi2FwU/Ldgn1CfgI5zhovbvZWO3vchjsbneKSJXk8HL1pIAn
7k1VGnqvsy7GkBuTyycWPuI4flBKZmJ65D9k8A2o36jhZvpMsvMY3DO/6q8i7hBHZ66pZRcdGB3a
hcei5lzRilNy9rEeGpB0XISNaSS7XPp/AwMilRFo9jPRm9BPO8ru8ypRcslUMurtYhOo2xSe8A8S
VSVTOxNy6RyUqM1mH0Ojo3mWjQwMB3BgA8hs0u9q/93rWRDEMvFDHHSTLqpkRQ/JjOdVfSYQUaev
PYdlQj2CB/zMywx0pNRQW3fQww+3aRcFLDOnTqf2PTGOzweKkR7pD+bysDYP7BC2m54BuYcYJdvx
x5iRCQ64i0v+AYme6ASQCzY+2EAeMrYX4IOIPgBQRMDc7uv+lhMNgB6bGmJpPIQv7E66EWa0QLHo
XDn48BttMf0f0k1WfsLqEQIdk0EvoqS5sXvy0tCxr9NhJvRw7+j4knlA2flJHKwjRt5e6vCwkOuP
sRZNTxRbYIjuxTDLfkLDRknsvZ6OQlf7qVns5pAxOUcOPyJrpl5s0ok5mFCCXksLWpr/jY8FyCSb
es7nxHmTV0XWw6H0LnAk71F0Bd+f1Fs0A6mVcw3An3XZd2qt855Tdg4hu8mPdyiZvqn0RtnVg2Xl
Q6ZfMZCDMpLN4R0f43enSb9iFIMJ+jaowZ5lMO4ThXbZrPHmBit6qgVfgW0Yd3Bw++P8oeCTssiA
5ayon4LNAdBckh9BV9XNvDB8Tj02rqqUXsQTvJdXpoXvWL9gwg7rjKEG45k17iBAkfJUVfvpGoE0
sW3Qduh56W+Qpg0YiehSpk3HvQnG/ZOOxEKa5910T6+CnhRLbSvXyAZGB4VFhnj5xa/IPMHrv3Id
XkGUaYi8OGL9Orj+1CZ1UbS9N5HzIz9g195E+oxGyida65JaqOOS4ZatK8lqt6z2O7z9V7uRxH1h
WeiSMkS645XAFEBgnE4mr2OwgfZ+lqASeYkK4vwAfRWDYlCncLlXhNb7aquieF34x+ySWMxLr5bU
0h+6RRC7VDJZ2Qgxni7VBe0f2LKFN9vQz4z4teqZ/cHRL6MEOYgZrdm8ZCkvrqYX87Ac4UFb1p9+
6+CpoFo28l/9H+udyFt6EzIhngwHHOo2U+jWjODCdXdnsUpXDEz4DoHuPg6ExAPPcsTQ3LfiDMK0
mnRBtlVH6fAYk7yVuQwWsFbOLuNv7g1xrIijXm3tCFwrLF3OhqqiIh7a3jHtOSIKhT579k1UX8Ue
chB+bBQBLkm04P5s6SNubV90K10Z7GgqQ3a3aIqRh0XL5U1B4Z4yyajHaAtLR2yl+U7PxD51ot8h
Uvn09ePjO3XzlISFLOConSo0onHxTHRCedIKCMp4/pMZxi7snIss9pb0bvYLbxdSu1NuYSxFSG3h
xnhhK5n5yqbmN+5vY0dUY4Ofj05IxkR7qda4FSAta+tc5ElMjzkz5O+yb9Ox+3FPPXcrq2L7uNzJ
DT3Wmw/Yr+1vQyPAPa6240CA2VehVSDb7C1Rmpgs8QaiJdp8tLoFw3OuE6q4VDR0spGe2lwgDzyX
sTN+NLs3uN4KJ5FcM+/PE5iBZUaqFSaGCmTIA8V+vzcSlrT7qH6qnCQ//4WJWkoSzLA/MKsSGwNy
fWxPbvX/fianRjCqglPPwigFN089FRC6mU2fSIe4SJarwU3QrRSvuLtfKK3E5NUUyCd5kfErsULl
dOi2lMWgdMJJoVcZb3GABW2kiF7p52LjKnBgHTgKp6dEeo4QDBiUGAXxoNqIp/eZzATCPF6jSv9p
zUAuvoovme+KEOJ1e4qFcVzUyffpPzScBpF7vpr3+lXSorAMFN1bb29i+vy0TRufILRLd2CbLaOH
7LB6G9MXiEYx5gAgIPpN/Zw+ZnZTBi350TLg0Zxm4aS+1ANCJDkd9VhImpQuYT5D2C2R3mVStP58
fQOE9VGbZbTly+w8pxe5NP6ruWflV3VVqzqnYWKKz3Jzvy4B/qBYWyvZ5aNYRYmzpyCFfUSTByVA
tx3OzRiKwo0or+YxO6o2Lir8L6O4DNFqaTRWqyditxZ40B/lvAl+7biaq+iBwvMgeg5wtMJlCDgv
OnH3zBFfcJvVipQ+hJkTN6C3DbT02Gw0yeVTyIby1ZdQKSyJVxg1SzQfZ6rfwJv55NHHMzt+cch8
e+FYQqAeRGYqF15rR9KHXvI5wBrabpafKQtIdVHtGVafvoeDH/U3eOGKtFYLnnZxhSKPdUxTWPCS
fKcDzHEWKT5P1nSfq9qkwSs+M4mfFbfcrUlrgtMdnaFV6npqNVgx1Hj5yZChgvVexhpYK6SbZM9C
qjmRdaDBdQ56bds4Z3mpPKiZVwiYoD5Ye3IBbFUMT2yRM9seLc9WuIPPWNzQ9bocACszfBAjAmwR
rpjeVD+KpDxSSWmpHveV7rZ7wYhRrvNvB/bW9Ux/fdbSecwYjlTINOxoc73BV3/T/sehA35PIrlE
OmzCV/48jvUGU/EIrWnp7yTdc1yLUwFfUcubxLLFOBJAoPx/FA4omq9KLTjwl04GZ/yAD6BJlXLG
Dg9DW3WgCBywjK1rLYCIL3vfDX4jDp70lTVQhr8IFeYs3GIIh66LebdUO3YWhqHmY6AdVzN1xo2E
43UiYN0T1Uy3eC9kFhqLwUR1XdeAop0XJEVUM/E5elsVrCU5i6WlY9zEElVyZJrWSSt/wOM24cmG
d0ggiBtt4r2n/MJwEVK96jwgWBwkKLbMERdkyhGVr39qcxwgJB4/svsIYCAoZZyIBCAR4rDD4NSR
d35L+9cdHEIvEgxgCg4U7ZB5XmaJBnS1b0wxZqp1Qf0ExwNDNkLsr4/bKrG2gexnSj22g/jORRH5
/6BnN+HyVnOoWNK+THv1JxTrnisIwzc9kx7FUE6kve8Wax4xjyvsRppyNdTjA2JZ5xYf4JsN2KIc
j0uQ3K5+FCbWouJOmebqD1QnTUvR/7a404nzxqVYtLoP9Ebvv5+P0Hz48fbBS9rQAlShvfkoVk/j
z3iyg0Nagg9kj2Igcvnw/guDVQYY321/FOf++7FWmyByDDdPAKAr/tOZyGSnrr01owF9iHwROePe
fBuw92Y2y8/KfH45vEPSAeyeCFCxyPK47HLl4beShqPrS+s+YR3WOeBk6R5rb3H+5OWKRDT2Wm6C
kHkL9OJMp6puv/1sOjRhcESjDbdZVddYP4t7CPoKFB4yvSUN8TfNfQ5XjW3o48svH4gSUA6xFXBh
lLS7f/CoW4a72CYuQbibhVs/BpuRjUZ07YLnMM9zxtzN5Qlz3jY3cotbdMZecNqz9zGGoUZa0Ebd
CfimSatc+lGLKOMdKXNlxqHckg/KXzZkdMxknTpRe2vZhaAlph6X68zN36eUI1A+5W3DOW7E6ywv
mPj/aCPOiNlCp69PM7Be8UekyrX3eBYTMdn8ekFVbUPop8qz3oPB6AWx4Sx9rrgyrcQYS4c8k0bE
pm5DqEsp4sRoPh5lLd7f+24EBYdpEWjw66JaHM/WzGBCYXnF4BPRFYOWZYwONxw8tL0xvW4r+8e9
SehlNI6c5UxDcgpfC+QwD+mL3QZw4GmFV/tiXzhm3CMdWFR2CN44hS7SOn9eXyCuG+0Or+WGeO9n
MpyG38Wcv5vjRp+n2IIgtlDeaPDDy3MQoJErFbd7XpUD7Ijc1U/JIRqBGK9eJ2E5ccmAUgleUApJ
4UVopBtdm/elDdn0eEdbwjGTFd9lH7ljYeOSDnFcV7jyl7RHQ9/N7+8Uqbq2WAoBHhp9mBE/dPBQ
BfGBE65S/Q426o8ClmXcyAu1qUaH/yVSwiosPHpJ2ImRBB8FWk9sQDOzwuq2JH1OxaxoyKBAsdht
NjFRGOfhwwpwO+G9MmWYOE+46ATd3yjnYbeVNcWRqLCcyBNCrikzfMUPlwe7JwOUL49jDfOsdE68
DT4bLTSXzeUaUcdLdXRli837FaLs81XdSmJACyZPkxgeCplmjaf74tkpnQon4hm6N3BuRDUJ2Kld
8uLeSPsYOrDi0/+Gnogj1Piwnfze7g6W2qlkbqVTIslh0oYWSc5krNlRLR2beqf91xRr5chP1C1l
Ztrb5G5dNu1UIK93WAuC5j/AbbhnQlvbIRJ49YW1w5PRxkvKjmapn+LtbN1RAAU+h059IwH66sHY
Rkd2+1hYfMUfv2BBpx8ahHOv5ecbhMIYiXabue8z50PgYAFMEgL0b9O8jp0BMq6el75atQzZ6cdL
N//Wu6fuKLNYqsFqHLKaE9enMpNDhfA6e/GNGVw3BdJdQ+mov8S7DIK/a1fUKcyNojfZ40OSPFKL
ttPjz6YYVRjuy88KzUS73INDgevUYmwZeatNo9u1LH02x1C9Atx99IXzC1E6NsmYjFkw/6mex1kT
yPTkXWoLLJBo7FNkLszFLXBTHyy7w5OrrcUHtQnLI3+F3i5CYyctz9Vv8awLYNvKR0zbxqZRcGV2
9nOCepiF8gi4yPb1HmCXxQKQmgiYpv8A4kUkGvXTawBLylcKW/odKcMPbvITEOiff0IPjSCyJSAa
JPSRTCrA2MWXxNvnWt4Xe9BFcThPmYAGWcLagLf8qL53YlWUCSZ6Oro1+CNYlUqXiz72ngzma/am
S8xRs3AGE1G8l43HbqePAGbLgN1JM7AvFw3qZlClWBf7z9DcXKGYAx8U27kJoLB+VMqFB/kTDTip
WKRZCm5IxHfV/+TeoDFJzQdX91MIxSLWwo8OrEp65aXUtReKMxiAz6XqAcKKwB2CFdnqhpjXr11c
Nn3vFkfSvHD/ZGJ01KoCvCJ8e0hWMGknQtBhmU9Jg4KQxPXD9N4Sl1HvaVOuqUaRJWkGlQIw9EwZ
klJ7xgsTD0q2MKu3EGvy9KZsgOljaJkYDOkO4ozF2JbeNHgzofL50q1EfzqBfxsAyyuAKNUXvp5r
WRxakqAfWgUfd2iTi33s6BQJY5BLjPTvBKc1uEc/SLhf4qtawvft17Se4Xc0jz4QgFhZ6QFn0sz0
l+XgTv/qACdQPoPXbbi7g8HUgIAPbtgcd5gO00TOgtv6mK0ActI5Km2MqZhJ/pIE9BWdSPCyTBlK
H0bdzE9sgexVFm1x9Iry9nQfLb73IWzcYyQx1+VTnA+xnPvFFYxMlB3bSXC5rMtIUu/T9MBjIrtE
uxo7qO4Y09Fd3q+vENzA0vLG4WLKoj76Z4nB+v5ru065Ontt4NQhafjsYtThDjLOkze5+U49dVOc
ZxirrLtDwYRFLG4qZllQSFatvtjDoeV3iwK2JHAv819RZV35GnrLfpTk1onmG8mpKox16mWsVztE
vNvuR4/w/19S3JWduREVe7Pg5osBXuLPz6JKRncLzxG+8vHBT2CEUf+8bcnH6yD7XxmWW3tcClwj
qL0jkfeWCx6m4Cy3xjbbg6FBDD+ME7iTQ8IVaE29G3XVi0SQ7lfZ9Xamm9pceJYUmyDQJDAiHe/Y
S/ebqoYDFj9mwAxxv8EGaWCBM5I4JQIcgzLrLmKoLrROm01b9ObMdC3lA+G/SNCZ2ycDP/TfQoUT
yAZF6dubvJMdCxBk/un/kJKRfJJe7d0p3KPIqk4yVCWELuk90/uqc4cXz+tXirCGppcV2x6U1ujN
NiFNb+TUxFsoOQtYXeUh4to0PuwEkseXrX4d/rkcKPZKQjgTytZSITsCaY9lPaLGMvB1IZ8EdKZW
MnlSHY2POZPrG5nJxHeV0XUP7CaV+E+sPRIVSbQWInuHut1LCGOC0EZE7zt60v6bU8MQBKB2FkaB
YI+9mSYKXpgn8kqVyq9kHkTvQ9HyhQFsrlJdVIKEmm+mXPAJqv3+KNT5QH0H9JpUW3QgXHfwAyoQ
9DgTt+dvMZLyCRIluRBnd9Prqz/0/j7Mvr7Qm1A/3W9aIrY8Ph4t9dPQ3mU7lI9mtphhGniMuBGp
8blU1ta16C1JpAyr8cyMo5Z0uYjLV9LdceNm+BexedCntqVvafo5Flyw9HPqMBdrSr+BWEQit3cH
sprzPXmfaIVEc8rtoXEEW7oAYDMpm2sY7a4dIKgLtwTBMyNBEXi+nGln46Kn+oN5PzzQVkzsQHkE
3FZF9GxoT7S6Xm8HYTwtxq0EDXimWdzvh0cxcSia8m/UR714xqn+M7ly+XWd4l6yvKycJRspP6Dv
CtMlByhUx1xrlLPEKrKovOjBl147i95k/U6zCWGCBkOSqblTqSwZCy60yy5Pf8sUit07K2jKESYl
m/HIlwr2sqMMmSIJQm1NsP5k9qAY4g4VO46/NjB8pQZHdtRIJXiNrXwhSIEMGhyoyljOcz0+tvst
TcIfX1i1/QmTsNaVjwpWFgtpzqXbMaHJj6DUHlqXCnEskqHyAHf8UYrzpghGCvyCgvQk9E/O/aRb
DZr7ozt0uVbUsFActkg0GeY3YB+mkvQlzcTY2oRC7Ewt5/5ZVutsebQ5c5uKyypDxShPTPI0z7Jq
myCnFemcvw7MCAgrAnaOCsGcgiC8ObDib0RDhSODP5BoQKHs57Zx7dNyP39gyU/TvdGj7/+aq53e
gsdV9rtyXy/OEVwnsJRvymgyHzGzWQBAHL+NxMrNCGHTlg1CeeGVIyeFhkBci/+Q01YjpOKUqcjI
rP3+CciDwNyDh7jfPvbnYhTCafI14IiSib3UEczmaUt2veEwcl6RImiZHqYRjS8Y1HmeTebYByX3
j3iaznkKRDku1uNzcRECSNqzXMWAWnUBpGoRmyammYqwnU8GXzntn1FqVCBiR2BJomOpqrmh/mac
5Oja9DuTTq26uy3tDk4aCjwxALsj3qM5s1LRaVdupdh9cW4fIOGZ2ozLBouFmrES45rjR3l7mWvw
BZbKqlPuAPIeXpCnzXf83K5L41xsYUwf6Q52Dmsf8fxVKrW5uC77X8bKMKyv28DWAFTbqc46H7e2
NE5xqh1rquHnixtgOB/i7fYZ8ru0rGaD8MHdPuwIxXVEdaHcgcdbO4fPI5Q9CaI9yL1/5PQbjsQK
SZ47JiUhf6NLZjBErUwLYrQdJv3EHEiNlWgE5TP/2uxwsrQhPxihkQY1hbepiOG1LfEdLfehoy6O
lGGw2zf+IAKu36OXmv9Im/mLmHEPA69EcYFuKZMK+hqvqmw3OyfR5HHWt3TGH+HoJr3yeANxcvKH
4WXpLXUzTQ11Rpjq+kJ2d9vEV4yj8rQdJ+45Q5qiSs/u/twu/5kGI0fRM1yCD/LZs7GOorvJMmO8
vfOuWiAeDlemi1ib/4ycjWxY1VHKhtcXYqf2YyUsGdodhUdl6Dt+96chFY2e8yAzS1e6QhE9gBHg
iK5CwChh5XYsxIVNoNsS0wiTpVlwjLvdguYDaGiMW4i1Xbh/F/9u7ONyfy1VhlkVc/w0yf+qY9T0
rG5JZuzeBLBMQoIRUh09BEsf8sMdbdMSqRxN9c6i5b4IQvDnaTeAPCJXUbJ3/6CnLJ+s4LL177aQ
b8ckNuUhMqMkdiWzjTabgerxMX9C4DRthdSXUdACtjAB2iBS7IVffQqUYXBCTqOy5W2e/CmNbYjN
wm9R708A/tUJnjaIjYDRHTqEmRFpaBzX8mczYbQt73bxXOGECRR7oXfbjpQbTVi88byVBm4TjrYk
h0TGyazVWH+ZUDEimryjHCa+bFmslObSlattPCohTDZi7jpurbyHGTgiOTWyS01TIBLbwy/m3I2j
nFWS47eUeKXCtb27ZEyXq5znzITeIN5JUj7KGGKOIjvw6FGlzHCJPwLWN0gH34CFE4oGRv4GUZLD
n0ksTuaSEgBPbUCMffxiLlTFZ9mwyiXNnEVBOVTQwGYwHJxYux1rsfaw64razmiCwUWi48aQIJ+7
rz5zuuJn1F3XBF90NBmmRlm+7PFC201FtdvW1A17smMZ1Ko+ybZNFoqo6la4A4QL64w4L9KvI/NS
joiS3vCgEFeBx142Iq6DDADxt816IXxBpFd3m7MW/ulh/SGrdQj0ntTMikZU6A/4egwvZ1c4mh0/
QmWTPpJ2iZgbH9rYwDhYmFWz3GIkY1FdQngtCEANwvXDM16quHZnSAWCVXnefXdGI7NOXk4JHSNo
+aAGG+OH7j66umuJmpkfL4m82ok2N/ivUhy+VbPKBe9PPHNV3uZZGzSQOKyhTyqIvN1cK1Ek0dXn
jnSvR6yXF405d5kbMm8jJWpFhpLiFOnYGPzHLDuX2uIaAqJsPR/wfuGLbgGtUzjkxEpILkz+TFwH
wT6auzAdSCaYeJHWityetH0N3DWWxqxYHbpDhQLqfK+YWRh9eDT9gokTg6N73BFQPHznX5l7dnJS
tnAyIInl4dqIWp0D0sk9DU4frLEC5MNqzvYbVGwOsXQEKi9rz6mLZbakerijQbcuodX15rKP3D9I
m/KGV2d3xJ8j/unpkz6490WLboYHjtxqrD+9JFFAvaxZQbMaWI80iC5KYE3Wa38MWzoMcp1DmsrT
R3gUX7O3/P80YFUWF0CkJvfl4aCkMRPEMJmwTdj1PvSyU/FtzeSFPFrAhUwYs6uLPpkKCt1iZyli
OhD7lPKqgx5GpXK2YZRxUDRO+Cn8senpztz7qO/WMpEJeZWmc51Km9mvZSo6bBcFpSFoxEPc8h3f
MDQkYdulFDvRAtfIxGiADWZWVVeW1d5ZMUPcpke8ot0pZTFrtD8e42wt0myrwuvMPa4Jwc2DqCyf
Xaln6PKurgHWkKGXkHcYcTe65Dp6YDsUJUXW3+hsr4RlMYGjrN4UXF4bkKDRxfJIhdkwwyi/QOnW
n5HkvFnmmj8ffUb8hmwFlmNpK2b0kQC7M+8ened9aCJkbolj3ceaeHdz/jCN5hdkY3VRR9JnqJRt
fg6nAh7Anba+rtM0QGaPu4KrdQo4wbu3fiOh3dX1LTMnNHxhF23KfbceTkgSGEywgJmE2jZ6b9W2
uGIQnofr29WmZ5yVbTgOFAcdozm/b2tiQ16MsVD6ktHO5wLKQTakTij9ztpp0xmJ1fuD067Vlpwm
1oKkMmZvPut4i6upDQEZcS6seAtbo0fE2LvGEAYa6tph/Uw6O0OVXVsLFKizOmzaUNoASSEG+3LY
QWaUfeVrjQEL50Y9g8Rzhaygro65fWPMVCHYJtTyhk4mvXo06b4N1EMmMFiGO98XTbaoAYXPglnl
KGpga1sEiFPcz8HwQ4wMw8SyADSz6dP/QKJelZCrweEqreWhjUC2sou9n38mNVW+9jsEymrqFGO6
NW6VJYagIgV0cEmboqzPU1x7zFqXKPfDO5fbJAmU0sWBzf/ow/BKq67zqf1CYlUSa9Ol4xZHo/y9
Z0Z7SC6vRmn1ZyUeyN8eQjId/z94YLWkMoDc0ygRE6zImAG1jllQfxgNQig5N4sMoDsDretg+R4c
+GDz+2+OCmh1gWmylViUGHyBZ4zni16gEr8fNBllndVFrr3L/OXOSykN+EEVlyUicovAgRWJLZGR
drRX5lYdFKLo9cFof4d+dxUP13gU3Xmfy7TJiPvWHUtEuThGswcYzamDzLIMG54Qcs2pYGmAi2mf
qhc5KmjPp+IQWDOMHEK5WOEcjAJs1HSjQHGwv+FnbS29OczzMcxrfXkU9+dWUYlV+RMdhTsfN5n1
90Kf+75lY37PRqU8T1N97c57g3lnW7CpBONtrlNus4ZZwdGzWbKDSTzfpB0WgiiTbPeE/SJK7F0o
jEgkEcEAYb7BfcvFLV9H/KJMAvZI8RNWxm1FKnOo7cP/Q+2lq1/1uM8sHNFf1jemmphXMoQPe6Uw
Hr0oiEO0U37a+L4J5OW1cCuyRFOxHbz185C0sMax5+E4JBI8p0OdejLeDegPYJ0uc+exGiAxtgOd
kIR2C5jssv+QIOlbHYA/m+zm7FcFWcuBa1U8jG9rT85uLfyiyhOP/JaBYlLJ7tNB5x2l4me+MkNP
rkIOlyvy6QFeSgcVD5uv2B/dXqcQLuqmixZV6/gwtPmuX0e1xjHc+fByQDBrurAosYf16hOdrCsZ
9KPKTQf/ChWBTenJdIZnDm/MIBCnYdS+jG06E/vRKKCLAXCOGWIrpP0z2omytVHWUkC/03KmoORt
yiPpDTM0lYaZ5AKRlQZTYLGDPmgiJYw+/T7ALO0ldZEeLDYSsAqA5d3ZqbNwlfFx96/55o6zQ+aF
kCvPNl3cNXcu8oDIyRSdHHAaX9vyUJwO59WZClL15K0GFqjEXZainGigqHjc/4ez1C9z7dtE9OfJ
7zPxv97yzAx4uQiakQEFqeApwcL2sIMAsdFYnCTYTJL0BhNb8ax8UkCNv6d914J+2NacuDK9tajo
gEgd+j6Dy0tIYhtAz0u1UZ5Z+sEh0ZcXyxK7rFhbv5SeysUdMIcx7U9hmmXG70e0OUehR8n2IWe5
i/7XXeWsMkBFKP30nkVSBtppvnfleLvpM00IA5S8RQceZJPPRtaCt7DlTT4vxFFpdjwVirrRDMTn
w/ABbELQeFu0zRX6Zr+6qi0KJRTWi+JnkXhFfM+/txXU1odlu2dekVaHFg4ZUmGEjP0B4/gOHNnQ
4i/VX2xhz7bZSgh5pTbE0DAmQEBW3p2J4ptn3MKE7deN37UtE27VojEUPFM+wQUAmiYS7mGE8yu5
CRyhkU2xk6lrVBDL7vr9UvyU881nXZTlSuXMmyFMQMDpMftQrss8j4EHGDbGwumSsgfEnoQInsql
LOYwXgXKItGHQZH9rN6T8fQleNt+PnOpddDNCK8qU/glF3Ze2HKfqXGh0kA/V6QhMo4AorscpoYs
7sPIoNorCNbi27mDLP71CZk/diHyWch3HJmSgvfgXYsxkHggeSUPDCensxUuCnbA8sw3aVilrEZn
MgJeJGUqrIzqs69gOoDjbOPiLXAuE2zRLIO3MjJmZY3JUbvvwlWpJbicroru/FJ/qO3KFEG2v5c4
p3D90JF3cHS6Jii2ji/4otDTZin+O5QhJGWRZBEClokt84y+wdtDYCYQa44QfZ5wzvpll1eVAZnq
ACBNV6a6aAQsLE2VKCD1YhG4/Z1dbaLgWygkI8IebhMn7QuAoIJyRVaDJ9kcFcKShpqRK+jt5hFK
w69jRo3tOkuggjJ2f1QvDyYWuGJ1tAowHtbZfi2gAClal6g/mhyXRbgNF6KVXUybXzHoAI+MWjZF
hxenup8qyA1oyeZI1ySTifLiyotqli6bSRuy6Ao6WpTZtF4oe50CjfU2ySOTHL2vYxtzMHbboquR
iLLWkRxCQNaCzJnKuGJMOUSPHSNmCRJAXfEhdVgI19g//BWNkJs4Hm5a3uyfdYpihe7WspWv7atJ
afPCrBiElDgsR7Xvn5idyw0iyeHPT5mF9A51nkLa+ufjyVkUQcSgjAhXWNyTC8OyrEj7lmQM0IHk
E0fyIKD/A7ZgjlA6l7E+IIrgos3HrNDX5fouWfaX7yMkBmAUFN6O+NDWe7BZOcvOIJD6+N26B7qB
A/0ffZNnoBKQr/NC+cm8g7QH799+3jJiaWzzUlc/XhJRUS2JSaUQAGpyvsDndjhOaz2ilg5rHLK2
Qaw+Re4AzMkovmWhQKSS35sE3enU05rmaSBsSLpcWhUL2kJRULcTBA4zL+56EwVKoCJ1/JJfHeNL
kXD7xEUvTHhKWtCD2BAQ4QjGuSf1Qey6QTkqmR8U3JfqlN+BuTqie3FwXXhF9DdaL9oWs9Drm1wG
A9kJ4ZyqEGPlWl+5K4LKP/3HQvWbh++zrorpAxqvkZL5pLlEs9pMwAFtjuYudAsxDVvLzFNhuHYJ
CEU9isPWObBYl/Vrp4WiFD2Kx42xYaQgbKXB2bvWgyyPFDYL7GVLY50R2yUPrr+BsS4CEfGqIiNq
cTtz/+iCvtFD0F0dQM011k/khYF1vHEcwK2iwleGiXWhOngfiI1v7GP1295I+UPT/WEtdpNA+25m
Dyf6otWb7J9bFc7U95nmV/2G2snh9Tnlq5ztNpYy38N2bt4sxOi5yKX0yMns/My3piTGdn7eb2yW
xn8ZnEK9VGG+rGB3hQHkEEABZbZzV3cjBMsxo11r2sHVV0/wDf3nnm8fgdasnpuWYsaXsKi9/l0w
RKJHfM9IQsXWZcco2HoAfMtOPZpejtGJxpWf53IoKZp7SO+bZy0Q5MKk/ioIQgMnt5n/YzNQskOU
aH9pLXOsXcWTsnX0lewaYvPglbvBKfBJMdUICL7K7X1p9Jk4aSObRaIxX1r0KjN9KBsCHfehQVyC
7SXGASt4d05eialGF65Nidwxy77TbQ42Pf9/dpx9l9nK6DbpFPWExRsBaSmJQuDfG5rfZZfvy+bH
UYqj+hxm0U72sN7I6rntJdmKg1IOwJzRG2C0nbaJUUKMPVUzfLW/2miQviC/R8WXn7Z/FtBNN8ad
WKK8IAET41ea/KFFDMU43U/kJX7v6EVyGdIxY8cgpANg5OgdAeyNAi/oi4Ur8y2pKE0LqkDLOQYr
Bjo/yL2TGZyTQRGMw4iI3lE2J4eoRcvVgNhlX1yasjNlRW8ZLAF7JRpNRdSoAAMshXj61Jvu6Lmy
P4krViUBBanRdbPIZIQQke2+tsHmujwaLoVW5JWpMlHrQVA4aQ/sfFFs9O8NJDar+M0O8I3W0I6f
4Bw+QMTGgaDZndezLhfWQ+MqNRQVUz1yAnRoYPwCiAatrQB7Z7ECrE4B6iLgzlOma4j/AtWQy4lo
BfVTmqnIJh5oOwUHlQ+tKy6CH6uWgZW/pf2eWTGDpd5H9Hefmi1cyHPxYA6RkIm6dAxI7efqbSN+
5LCSR0Mfm7SAFtBEo17rXxTmNIFpJp9Hr0JbSAYk56+ZYvfbFFlAvHXEb2WlTFJ0sEQ1dHy1KW0J
ew/Mgbs+lv8gAxv7dG5uoIY6Q7WReaYsV6obB9MJ9jO2RbkKfpD3RkJYCT6Am088VL2BlNjHVX18
ruMg7IskKwnnmGgjmb03Wxe/fRK4n9WoG6F0gCeD2/Ij9ICRY401qFn26qpxruViONyEe9dXCGSf
K9SYB9lP76x4I/St8mcOm7QFQ/5M1lbrcHu9Md8n/9DBTD+MC3sfHVxiNw7BUXGx6F1G9N4UjDE9
ifwZ1PxAZy843ZjqWCepFz618Q1wc/2O4j2nyFNu+kvpvAgJfD3pBgOzC0T+LvWKJARA3Iq9G8I2
AkBA1wwje4fojZD6FLrkQRUNUtzjXb/nmevHYQwfLNBH/5wHbFCEnN1COdmZXOOxj49Kvsj94s3J
aELMtQATr522WhlVJwCzqYInItFwmxqelsTs1bGA9lBFPpUQMFPDvuDofwZtnjoDluLAV76w5BQL
bbaaW/MROouZ8az1msZAfGTA/Bw4njYKxb6Gt1a0RQIrBvSsTufzhlD14lWjMstCvoN/QuLC45B7
hk7HI5UxuAaDhb63FJvcUb7IGCovx5BJLRJ87KaRR3MbYtBnGbD3eNtDvViq+HKRGOXxDJCyG0mq
WFEgPudyai331XHFnkNm+/8IP74B/n7ybdDa3k5rKNMa1B68py0xJHchBWd+pRklOjvn0bdbcgEQ
0+u7r0ZAYmyQLz7Fbe0CKcrNcOgqEcr+/z5aqijyhYwwYld02nvNVzHhDPE+qYPWEotZwI2RoQcy
8Plfm6bPzY7K5eWj1yElgC9iXaP6r4kzfEYYH2fjbsUERc5xLGCZ6fb6PbIiXjRwhvLoo2uZZN72
MXSSHxok1SThNT/w07Q+bUl/OJl2QrHubded/p6e5HRki3Faly1i5H+6G1nJ4jF7KFcY2oaVGak3
UglF8T9DvZVf1ZeITBrJt3ze6YyAxVUnHsjwjxIElWlozvAO5kT61WwXOCL3oKt+VRRG6kv3RZKl
FTR2J+qg5uzuCUhxMYtK/FvGboGsbTsrcZtJSwNsuqEGERiecWA9EG79l3IokXM0icT1IZ/XNHmt
ciJjdgaicaIa6xqIKH7ywiqAZ1bGtFuOpniaJ+midmHb5DBc23gVNy7fXstkseE1nxpAPOFfkJgW
uMJ7A6bN75lfHj8aYI2h2ojFodRG3NItUdLgxsKGflP50jWDLHbWHKSRgysvm2jYuEKS+mg5XVdX
uFoSRpl5GM/ZpmeD0wR4R7szaoCRyVjtFG7qExIOMSOc2FJKdmbi7WMUr1ShYTK8js5RIJ+zeEwx
gMZN/ipvOLuqGmZUILd9wNTKhy/veqN4WpIIreRMGMjq3uNMnmVnECIEPr75YrIy3TSdrMbV8bzd
XU2FNsrRoJVGpXtpM3IBDP8WxTatati9sRsa5VHSWi7IwaYrmfnZkasCPmnVyKoxjOMUj1I9a/ut
QuAu01oDMdXMyXQY+SpMkizFP2rb2/J7ntPOoPSZkisVGGx3C9HaL8372J/3NE9QosKGvUSwygvr
Y0gQbYuwKKwTubAa7bKTy3Z5gEBPUupQXzzeDnx7Bp9uqTm7cSMYx12mAqRLl69jlWw1No8beYIp
J6m93kIktQbv92g9J2MgBQiQEjM/1cCYi6P/Eus/45PQN+wFX7ICOIlf6WqLoXO+IuKhHVvqkvov
RVu8UHtumiUbSCdrGhaAA5RwHzbP+g5jN2C3kykq7q3wb/Z+1dyL6cN80BQ8CzAjoKS80Ac5tHMg
TmEFqYFJA2g20SjyEXwzYsgK/c5VfbG3KFNSm4Ur1+FWNZG7/7p39u/9y5HJ4Nx9cwwE+RzCQqiK
ycgcpOwSh7Eb4gcsavU8nv5LDGei1hEH/KR7CrBEIXn8xvvniwdovEmVTR2hhKbJkEWLq4h+qLii
SJ5cuayQmy1A77GiX+ogqBTjbuWN08Ub2htSrsUbDjE536DmqnoHfLU+JXNsD1SPy3Xex7usycgf
36zNTM+Jo/fnUggTMdBxydM5/MYD3RIKK7whVZ3l8DYpP+qWaEmMHGjaxeeGVP1ahpH9Qrz3Z4V4
0Ylj9NxUEqCETorM/stgCUAR/KduCg22akXGfhZbrCzOFwajV/BZSnmXlvh146zdPm3YPQk2aFkX
LxB/7w7KHaM5jQ0j1c6faburpkeuLXVLqTdy/vjaNCBtwLlfSYg28GKHT92vyAvT0NEL0RmqkYum
sHeWB75ZBi6Jh61xy//+k7ICCg0p1imuMOjZWNF09EMjmn32HxXH7MQy1FsNTlvVB+O+Me3eDiDx
mT0Wytbk78YKK8PPUQy2FbdHycqca1q4mi3Xx5+5uGIiKLzTWS+UWa9zGNJsvL2uBkmL+dVRLJGs
vO+5nxG2aCxkDULTxdOkrA0OV4MzWslx2xl/aXPUsbZC3G7XJkqeFE+faL4kfkZocggX+IZoGys+
exhKvvEWsb8dUaDufT6eHe56LLHU/2njOEF0RrHwYnXpgRwgRDFx3pSHyZcGISgUiB1cuklLXys4
ZSqJ2XLhzl4lqh0y2A8xLatY0TDoJSATXMdhcE508S0B5XmAUA1JUyYUe3UdPD2ld0qEYDDoyKr6
NgLRNvby3mRzmXCV2dWodj6pap+jBpoDsE93WTgLTgeCzto/fb7+so/fSNeNxaD1dylJvNmenPyX
DmoZJTOoAQeAEMv3o+diG93ra3XU5U+8tdcNf2buDPPg6jQEMPI+KiFE/hWVR76598CJDQoAb/+T
1W7u81wbZoJyTPJ0A7NkTax4mKQIZvb80nZkI+dRCdVyvH3xcG0bGa+XNSN/Goqf8lPFDdl48DDr
xEVbEe2AZFd0BByiTuNO0JyzBSSDSwT0/S2uC78jbMjWx7L6nErFstcqb1Gx8NNoJ02e9fa25rde
aa5wyH/toydrBIVgzpWaoLZk8cHDcLkulMPw/iN5bcgr1evcvAf4bV7u7LRnU4V3QmE4k6WTi92p
Zr8jVV7njmoddhxvg971va9Bg+mqJ69yuT1nlGGuRbuD063Sdunk5rmFrLF6op8m1LZaO4P77zlT
4ZjisUQ/DCUXjpZtimoshlzwnTtb7W+OGlXF3JamvkNqBI69Tn80Q4EDuH66PE3jFRhmc/OpWagx
muiN64jakA/GC1t5tpqekLrnJDJW1u3zFt4qjIgJ90fWc2uM4P8xs6PMDqsTriHTPKOd4sh0t8wt
QhZcmVhWdpX6Vll6Vp29o3QeHWgun7qF0ALYI+fcKzbSN3HPyVYu+b7lzZxDPb6yjb7MuZFbusD0
2k4qjWd2OZ/tOpSxH0J8bGoJa4oT9oobY88XAm/PGkJcra8oNjNbWyQQnNwknyo/oA5uu+uU/m03
1wr84hh3foUAQTiH+LQrCFsFvXL3256GLUu8bCidb/p2yYELmHd3S6AZzt9qKCSOYEzhnVPdJjMd
aOKfLruUgo++7oZnmbbwq9Kuyr+R+NpL3gj4u1xcHfrXMXaN3Lt/3n677E3zQiM5I2Kna9A6LkwY
7yfa2xRZWj1GpCussmZ3Au3XkEwiqssGz5y0rOGTbBcwh1nne4fvzSbikqpseyzRjQHEmwRaoElH
gf50gYdCfRvm8hizc+ImncttmFWyWTUdCW7XzWK548yP9FrxS5O2eKYw7Kzn2so6ZH8SKvPH14PO
wi+TBqSanku/vs6UseDv9l/xH1a5MvOFnx4ruUZl9XgPVw/eC1gxSoFDWOEZhNtsAG+ZUU97C0Ds
odpDjqfa7l5ydkVGSJxeOH/i0dTzJjRUMS6r8J9YXj7CvBW50ZY4kOYCkM/y3VduVhjjHCLbIqMW
v0pl3gKz2y2P0arkqwlXptGjLZTsoJqJo7oueTmQIfYswi30MgJ7JR2z+XNu8iqvG3SOy/lg7Qnj
8EG5j+lqJSiFSh98OG0RFyo3QHFOEgshSi4oM215S6SFkOVTzI7Cl6rzwhxsl1pmZxzsEClSi0Ul
P5ee30lzkfSMSYwlBTAyvllbIMD73FsagYN7rAKM0ny9K59Ij5Ju+sYkEXFEQ/PI7s53jXDr506n
RNMweJfyHdAs8EZq1dlzU15Jlp4kTA9zrgJzavRWPPXgYZAqTF0DY6cP/rdyQMehgDA/kAI4ZDj0
qXIBJIkZ5Cu9wneaoNSEcTgZ47u+nIgdIHh9NkCKJq8SuPTEuZ/MpFFd1WRhw7Zlg7SZM+lQOhkl
9l3SzHYlezcCdwrsig36sv/Mnwdz63nSv5Xp3lWtMuV5zZX8NWL+4IsGkZdUTLAuWHZYR/IH0co3
a1EZl3uDS8BmI4tcvQL2tOCNBmQDG/uTQ8INyq/jrEBAZWlZDROiPBvVSNlcgfc3uNX6kOAzOycv
llirb79vPU15vQqYaRJuXl/smHy5RynY2Yl19TQL/5QoTfDrj/3R+uXEvx9HCfaytkAcKPb5Wm5s
J3EqIkOKnm1rRUZ8gCqDGEVXbWW1qflTo2BeHgJ9luEmR5EkvuijKWxe4n06/3QkJkvfqY2txbxz
oUIQnoR8O17JYC6Sq0AlNzGHlPqr8MVyPfCqmHtlqGZ86AUAn+DMGFEFPhHidEsV9xIy/OK8BBMn
4dt3PJWKkrGvZuh5IM0PlQA4JVO7SGZvi3hrI5h2pCGt9ec00E2vck5Oc/qW4OpDjH5DtI4pWrRh
3y6MadjmhnmxTPw7M+IG7ukvSqEBAgkrU97gEIN0uY2oz9IbltY883vBS3YhUZl/RVjl2oLQXe1A
TXyfq/uqr5GJge/cqnecF6klrTGf1rvxyBY6hkaU+nV2cWnYu/PFTjH0NvDj2+tgXi0XSk8b8hq5
xOLkMD4eQ3HdcKKcZDt7e8ifjBf1yPA+PIgNxeMGDz/PEMZK/b3akJzvrNkq8HFor0TGRZXDf++x
SxKVjPTWNXmGTek/oiMT8FWUBmTWHXZ/oOj3mHwxDT5WXWbm6pZsQJOOyZLe4q8ZX7DHPbSTFHkn
ZwhVjZk9hCY/6rdtF1FXXJxZB4m33382g796MDp2I9AZsvRvB3n3DZzJVtjhX0jwRXabk8Fv+PX4
qLCT2DZD1AP/Ez1K/Lq/ed8GudKxYpvdiPHyZDu3lCwLjdHQnkalnyMGZExnSLYHLX9McOZEiq3q
2nVVSuysCH97lSCIXWg2oflLXaQQUHVFKS3I7/Mt5L9yqWlhXtiIdT9ceiCISuvJgcMqDDtpfng0
lPMRB7ZDcYhWTSlUk9WV2M8T/HYvcuX5Byxqwfoscx5AGh0eyPFZP9nqzw83OibBC9ylXbIaGhEh
vp0BYTrDTtkZYnp771GqZEfrbgbj5eA122jAEr622UsPbB7gv5rykCyIgD+ueflXXd96m3sctCpI
BLyXIi9KhJ9/9/7NyekYLVasMqaH+bUI39bS+rksOAAWV+3Hhc4vTNLSlpO8rrksRYc7c83KU4/c
hQgOrQYibuWIQoPYTveXtP9z3lq7u5cIDmlfvJ1o9IO+SJp78/U4ZdW+oLJnu218tfgqC9uIzJqw
5OI00+J7k0z3me1rxGqZI7pghhbaXYVjCbr7y/Pj7gc87UMBGK3fc2+03ATwVjiQaXBuX5lCyE5g
kMflxfwRwGSSlNVOl9dJ8TFl3SfmzX7Pnc793fc1BD9OvQbw8hkQIOJABvPky1BBiYqmSW6+Hjby
2gs2jiWexNHz0se8zDOm3yeTdal7rX+KlrhR7HCyxTSLAJMYrZACCp2F8O7ZC8FhOqsOrJJercZc
dqOvNMiubm8MnDImAON4Dr+0xWmBqdFRMM1JwdwpSN0PcHcbQQO23Obmk5PZ87+SExjv3Kb5mpqc
4HRJwIxHQj4rxdb5xkJSnO5nwVYmaVPW9oOhOaX0tZ4C5gEgPaJgJ7dWMffTqP+eZ7Ye5bpFZuq2
s0JdzucKC9GOZ2Z8HLFUj5PVFnemEd6PlxElABE4ih28NK8bsS7PB3UzZfagRWUKAW42Z7YAxaxI
uYLMZ/disE1mv14FGsb5G5Tz7kkiPyC4owNcHimIaFpNM00wR+XrOvIebVDRbYK2Uf0MvWKXajj3
X7DRqo8vbcK+Swfr8qvh6i/KEovANYxUSjsc4RHgGcwLTDqKxUY2zbzg0UXAbMTG9A5xfBZMyqcK
jwuHRPuXloO9s1RxVUM/3fJroY8FzXKBCiBjg+PSK5K85rf5+NKW066apoTGOY0xOr4+6nyWfFUx
UvofSX9txcFOd8Hyt0j9ZGLbSD3JIpfBXSgqWTbibOjAG5Kxm7kRIojFiuCtm+uZa8vH4/YxM1al
53LVTjmj1XcqhG3GtFFGw5VAexqjqZIhY1Spkg3nNyz6u/wMA83CuRrua+PJqJexV+52xkU5rLow
AQ1qKBsItuBmnYz5+dBEa66qUm5raB+ynliZL1ULtbeDb2RoJ5v4EP3sYOgNIm2JrKzkr4SxNgV0
vD8H4whxWF84PYyWZD3WU69sD+ZlCRNxxKsJWSgFaVNodZZFXjQMGhm0+eb0gA0XtJOQqfGsbcVY
fwL4p/bB5sNikRLWIYDh1tJbNtGRKpDArLc3HAIi4nxWI/y0BERS91Bsg3Jenz/D5L8JonKnPLTV
OHCcvndusW4AD3vSP1SOWbRr8VmQcB7MSGFz5bUTGHeAB9BMMxuEWRRGkbbJU5B4xFaoMzCQo1Ob
Fl+4AJe9fg6CTZ8tG8Lyfg7vR2Fzo6lYDIpdzAr/ogs6VwarLaRO19DyL/c/nJm2PejGdGFnvGZV
Yhjf0yUgCIT1JFvAq/cBK9mHNgEKCG7MCeMJr8TzL+ViJX65ImedR9WqXGmcPx5j09s+oxeKiOX+
l5GMe7Ol+ZPCVzMxLTOQl5bjiadhRdxjnIkz4SBFf3i0BJgW2vkvEEd7zK8NJwrmcJLdPqhF3+mB
bpdq1xRAGMewXqwrS+tGGskv4fslJL9avrezhVzR3yU5CXtNlagxpC/Z/q5etvQ9tVrteypU7oxG
qSo61CVMoFzqkrqUVilcQkwTNtxPyp8zWfTqAEB4gajxUGbQWtGgJIQoF5pt9skIiO1ryB2+zXe6
9mNlu+wfDO62G78tY0aGzBDKfle1V+DBFPKIPmpFsL/vDlGc74BiioADcg9pJCuaDiMLsFRkhtNu
bOPthA4/SLAtCs1qIQQbhPDlEYkcWxLOb9Tgeuv9KFYes4eLrxjSz91Z7a2Kt4W1ZRGAS8v2t2Eh
9hklPbVqHu5nJrUcYP9BCJAJYTg6KzsPucWGlISZpqezfbwfemwvITb14DDzQZay1bf5EoSfE2aB
Hrktk8AE/7UrROh55bz63YM/x2e2q2/mogtBD71PkG6cDg4Ob0HoeYwXq0DSzeCHb1bxZTV95wzT
dys/rFvHRrF9gPAe+oPV+4fKrU2DpVDh+crMdfX5EtebGW+va4VJVE41dwMu1Q0lOkmDBKQkz3CO
p63ysivrl47NNLKWxCc75YACRrpbSUskc5X5OOAQFZtzdzTjhzs6K7BDJ75fxY6Duwwzg8vH37iQ
08iO21TwZkfNzYqj4vNzVz274gY1/ZBBwZYx/MwjVuA2NE4JD4VCJnM0D+t3AJ7zvvdF2f9rs/bz
ilhlQfwQbp8j2rGHRKyud5ABd6cXBrtNHlAV1yfgqjRFtv9bBF+WgP5GV1Fw8UV/yM7frhTh7AaF
iJlfwBMCD9F+hblpym4Jg8cXvMV/x4RXRU3kS+6pDlkXM4QmBMOLcSS7P509cr5gIBeCOvOFzank
HEKiJ0ZX0arRp6QdBq/IbtyytE1RqYNY3kPWBDmVoZ8Ei8PqYQBuuOJTB8WAIaHzimymPJikgSTo
AkK2GPNlA3HZHT94ce/YVoTqeZMHsxkJvENP/tbbjXKnpNEYcQw8Ehqg7yXEp1kxZWRBkKGyszfy
4juSikb7Wr0s88/sB0LUOjLMR7IrqLKpZxCcg54jTOBsru2gSzYswMGhPIyTCYZTyqdetRo8+j9F
R5UdD4J3fuNd5gAsheyIy4weDAVVwvirFrd2/kWKdYacUQ5W8eI/3QuIX2i3wycC4iDM/NAij6sG
njyl3VKVvP0onvCnUmJwp40LSkx47mk33+AlyG7qetVVysauUyBxelE8CCz58Ut4oic4vHzPk/Ch
r52NnJunLiPaSJFl619ZMQIZ3I9xyIKlW13pjbw1FyU9paVGKI/XpmeBctCbgujNu8A6NKov8u+Q
sJ8xzGY+WaX7OeXmgXESI3BtKtMgPJApmShW87FyvkGxgM1GzaDBXdkJA4fN0WqK+lPlFY9kb7u1
OlpzQG+ltPOqKI7jCiATuU4tYqS90ZemOIWgv2z4Yc5d2i5HgE6ZW04CjOhJKdjkMqVDaA31gLAp
dbzwvp/EH4US5LRdlacdi7znO3dmZinQ8yZZvuF9+KhSe54np/SPWQTfe7cFQcTK5K7G8qJohOGa
bK6EwU3vjwU5wC2F8Q8JQTzg0WwbtHmRVUlyBeTLXNXUgbcSEDYMnFIRtrp5ZssUwMhP0fxQu2kC
0q+bTWw1a6O0f3xY8Pqwx5vcJaeh9QtIKuPRoHA4uxI7SXuouH5R/j9kwo0mAfr+SwQUUxab5cyt
siYljDGq2Wp1rwNXiJHaaVeA55+YEL6BqEyI6Q8JM9E67FzAp03kZtbLFxo1E/CYGFYM1K1DqRSp
2BrMZEuDXqRn3ADq9BFGDBTy9OzW3uf0UOPLq3PWApF0dsItVyZoo/BfI1hXZrf3jiHB1VEBauNO
wju4mRWoFejoV21c0QgmrAVuGJXg2EmdPmbjDHOIHWnXujbBugxdIW4FOf+EEN62Po0iXOT4ou/b
vJP9jCjPoSWLZiZzHnX4jJsuwjFFKjxENe66wJZ+SK33eq4mip9EBx5Cah6E3WTRqmkyBJD40oyW
TU4Hgi99KSLAaojTX+zEm8DucxwmdLJC7p7yEWRyNtwVBayPA0+PHbhGbOmIA/P/RojZof5egHvg
dYF/gXYUJsWcNeplUUyxisvvWomoMSsbvPbTmZYujzyM/zHeWlOcID+TAQeqoXinWQ+/mqsEx9MI
qfeqT3VXceM4oJWlhswu/8PND0SuFWOx13tE3LplOD7n4LuaaLZedmC9RLhA/IOkhThxOSOydwho
n3uvCjZQl5kqBCuhZN/L+KROzX3fVVJ8LaQuiDMM/g+HMN7IZquEqanhxYBIX7F+x87GN+KtJMa7
b4882Nb1BCBgkwGPahM9MFYJG0yi7g2AZQ9LAcu1x5cz5gNm+770bNWda55ASEengqX4aU6gfNGk
luBlSn0DIMs/COSJCxLsEyKzivYRJ+ozXhgpsTxXCVXqErHG6pavTNinc3moT8X1ZA4Fw48LlhX1
0VYxX5gpnhDi1GfrEVP/XUoK5JxvVu7me+LZYSGro1OYJ1s04os5LgxzixPWmByBy42jqET3qZ1u
Ms+aacJqFCyVFJveLy7WFqOaGvsk839bXbyMN8HDf84pMyUVlfEvh1LPLzyOwveZCBRlfwasjW4N
Q3Ww3w8McMjTCqJzB2Q/mA/yVKeeTMTAnotg6aAAaVewM2k2lvafrfuXfq0WH9enrT8pWksyaKGu
YDlM0prOz+tGoMaGVOqU2aEtjctbWXbrPklvaOmvb9XWyIbdHmCvH+lYqCAAKmSKaoiXYPT83PJe
FpVaFwcV9zhpgmBOJHu6x2eurWD3GdTimCNijuJRstZwAemaqcp+UuKVHTaFa+ZRQh1Xe/T5WVR+
tgCftggEtf02APJmOu6J87hUUsey+BMpQPzxF6WHD1hqs0zyTO0Kq7CLe1AiOZE7BnX/vuUtxveC
WDDp3A44QkMk68HEHpsThx9ruFrGS3sYLWYYXjVe+CGhzyNMjeVcAVqi9GmaByY90kuy6e/d4+sK
I3asBTDBI/uB+/UbtjEmEb1UhsFZ1xDa+OkkQKbHZ04cCO7b4Cf5JSqlxIi3cTMv53ftSxokLRzt
+KGkpyV/A6waajScDT4Q8BNUQPaFN/q+xfmu4n8H/qt8JU2PKEeATzMruV5EzRSBpWTLHOWXD/oi
I0TIsDcqqRC3Tb2zgCknMJPyTVCwimKGLmn5RgaNQSrczJz0s4rA+qdIfbz3i8ZVHucMZW2mV6fl
7FaOaOjxItPUzQjJLCfdqatyI2ssmxua/8NeW7p2tdaXQ3Q1sPLNi+hqbWE9+fLPpV2rwBgBSthJ
iJeTletEWm67hsEEDHB+BuraKA+DOgba5VbkAmzxVNqmA5brN9g1ZKSYL4qHxfCgUmUvGgjYFowM
PWEkHLT1BYO3pJFKBF9JZ/SZm9PuN/Yj/AwWYdM/5KGgEJzELU2sVdcaOidR6krTmsLm9wyQxVzR
3Qwj+bSTakn+sNr/EwNfBqVCV6nDHCWfnS6eME6frbFX9KF4TagJNi72dDAIZtggGxZvpT4sFaE5
th/5nZEsbA/jzpsXRQr3iGRHz6+LY1HZjk2MSI2BoWyfZvGFbnJ9exIstISZy6amSE7+okak/4NS
+Z13qkHrT2J7VIQFfptaoc4GYrBbL0VtGPeMpnkuNdEJTufMGUShZx39xOt9S/qokxT3mJllRnHP
LJIkzk0i72HKlZBp8kzz735oYH3oQDadtWc/khbHNDQpl/zlYeJR0vsEiPfUHfenohfSy9x8m3is
3kBXoCAPWBQFLT+yrZkdIAqaZetQ/TLCl6A5eMcgQqmXAAQ2BOAupqnD78EIdVjd0c5xgr/481PU
zAC/J7J9g8CWpgHSs2TJYK4NdRVkg0p2HT8CMsloVW7zdjJsEr3LtO1ZUwqeyYQ2WMnEW3Kbi5+X
oA1izC6JahJhETjrjNZ5FS+TEZ/jYbHB4CC/9wauLxamrmAsff4DPThUG4roXb0Ve1iqjP5YOHp9
+2S6qUs72CH6JM4BYyKMU94nly9g9SrNTzl9PQ8eDbNJt7I8qFhOVmoyEsqo1RKJM5DoeKuRrL6s
qfoU98xcE3a+01Qx31GbyHEHrXv5G6hAqjasSNlpQGt/NfzlVMo7KyLSlQnZOMMUBGfNF+jKzjzx
BR2rUUvkiS2AXVOxcBr3xmJP/0MEeuwy2IwpRFwpOg/Ygu1CnLd7M+A/9dtrbadjC88sQCp9zDYF
ui4E7qq+FD2TVOLabGqa2uRPO6I/FHvPYURGRz5Wsxh5JcRdnptwezWVL8nTXhmHPqfbVFhRNBFU
U08LNMkBfgi4Kny2Sr+nWI4YKCUAeHdK2MCrRsOIN246QxN22hYWXIthAqRl5XK5eNRlWeVGYJbJ
uZwU951n4D6Ouzn4QJaCKsfKjTa3WkrmN3YKp/TIinHBTP/ey4lLJ4Ykbm6EbOzzlMAW5lytCSQ1
P5ETQizxwAosMiYoazL2sgbJLQXvf422Jl1HWTAB/Kq+jAkTy30J7dtuDJPJUAP+W3PQKxbhNNPK
YytDljkmnmu53OQHkw18FKCz6QG5WaLgkIrVjMGsry3KYioqfDEd/VCFoRt5REo+X21w6AK+9zEg
igqlSp9sCys7ZiiFavZDCzWXRAd+vi+wmu2Fk+45+HyODwgAGno2LIWPgaRPX9Sq3cFq7eFp+T8p
LXmNCuyQ+yftLm/wNF6KQXSA4kfZBJdONxkCz5b701BicOGJ8QOFN94M1Urgh8gUgVqJ7/eYX5Da
DRYbUZsP3Cj3Hf666V0W9X0RRDRmVO5/1cceM1YMx/GLzroFHUJlQemKNBJ0suwSrrytwRdTd9vC
88ziUNOuKeycu4/TNV+iMHjyk9AFHEYrou5Ynr7cMXRNcl6R0GQu3q11eVVRx97bKKluBFuQPRg1
MumfPHVrSRnDVGtsCMQKCODBbjHtwcQOxWiazR9wCqA3WOli3V4TIpcqgxoC7EzBw8s/qPJZtjQd
ZohfgxyXPsb/f52w4cTtTMnprDQNZmMpKqHcwNXUdHHSo6+4/eSkGUC6YwJEncaXCrSXbp664dJG
gtrNQHs7mqclefIHTEm5dz/vSVjcyAZqIWztxkBjB1w/WYqSe2Gdemd6+Xv7RJ36nTVQTbiyFXHP
4CQFFOP0VTLawd5bsp2HYTAPxD1T4zkPQMBmX7zX/lOZlaMdI0BCzitpVi2mrrtdGbX+RKbJaUF5
M422aNKuhkUVdCdQxk2c20GlnMa2xKAlRIf1nRHDNQ1j5fmTpxGmaxIaupJ+Mf1Fei1WMRjDwKPS
GHSnl6Dt3bC1D6lAIFAoDiogpZL/r/ghWOHXPG14lhAi/L6kFy9ktadEis+oajJB3iGXiMi6/9u0
okBWfH6XFnfM496J8RViGSjafLuraXgyZu+LpxlKDzNZwSzTYd35Z828VVnMYZldAlYzGlMlECNc
gu9apxRVDxtSsxB7ANviA36QKYKiP6Kfyr2nvhW7ThoJsVbAE8GiqDzyqJg3MDdeV0mAydOAt1RM
fKcKj+HUQ5dCgbUxu2nA30ZCUFDEU2d1tjh8Ww1+RhpA2eyU8RG/UM07cRsiBE50TybHT1vKV3bO
HBS+3sxqcjBDUm8FPJt1QUiydvY6wfBMtl8HEVp3Ui7D3GqykJzBBq/ZUSyUFl/tAsfYSY4sy/3m
Tzp7nEOY1X6bKOZkOSchsJ5JooZ3PSE2Giyu9ol8UiEeWaA+SveO+yYHBKDYj2pJrfEbJN5F5EHs
0yKsjW+UAyHD4mOIFL+rntbzRj5OaI12WiF3zkeb1OTNJScZiI/0tqf37q9ZuCs+kEnttr+X7cLh
fJGgJteDioaciBKqBTXmGcr/5tWBzOAEIex9043Eg0gwozLSRJWF7O5CNA03BO4aRBmtkbO6NYnK
8q29lrsqrRLlBY28lBMhgoZnwYfjHygJ7WklAlP5n452Mt1iSZnaciok4dYNdGtFljgVNIdNb2uF
ngE9igFIItlL5Cu9NcW82gNxLrt2CFt7noskRPoQQR77R4Tfs4evH8MCbpxtzx4GaUdh1FALI28Q
xt4IxVbCL8zzHEIikQuOLz6ttD4MEH+V5wimq2wtUVuvULwTKHgHEQJ3xYoERPUjHGNKySzVvsvz
yNypSNw/n/Y0n8TigifCbKXjoKYCMXhi3rPwsIn0csHJ9Or092gi9H6sBH+TROfzQMe/VobCFGei
CZDD6KZvYAUZOnYaCFsr5kO4BIQumYj8FxZs1B3gSqn2ha8JEnt+s2aVozskI5bcypudoR3TzTHc
14SHAEAme50+5O4IRVPpk6ap0H4acF9IP4IYSA3ZLku5m3/3FBczoSlasd4KPDuZeuhp1KA2y7K2
vaCHf7PQ8MpZrd+D7Zas8zVZxUtEgC76NsFEmam9vz4TUv4HwWUpFwBD2SReOnxb6Fy66oUJ3j+0
PTuHKmuTbPwB4B+LtHJKFu5ulmHeg2ukalplSdl3/b8j5bt3TEn9HZI7C85VFxobKucFAaoOdr6F
dSimT+qHetUNi1ACsz2n1UvKT/j8DYmyQKbsxPUMeh6RQw+1SJ+uVP+PSiWZZ8sE7Y9+ZGWp7JKo
GgHzVyLckCjrR0CXqFMmmWxzIhh7l8q7v4H3Qiz+nJDPT66r9SdQ/mRe87xVAsHxu6WkVrBFpgWq
O7oUysH7WtF9npZ1mmo7ySDEi1U5SG6WcOgpIfz0DApG5VwVPkbtrr8yHjKNie1Tgy4vpt7WnGxo
5jHEwmcOCD25VMGKIWkp0eokFBIAuIrXJ6zdh0RuDwmBrLPvQY22LB7tYEK59wtPUIT+5KjLsaEc
fAivPzBkTl3W05PS14PP5Qs6A1M8iLkOSFUmp2kNY63Kljde4m4gwiqje1yJdLQSbF5g8YvTQwZB
9BAljSikoa+g1C4CUpJXXBti+6JTMdoK5rjk4I/Et9lLHhiJOcRN8lQMT508vjI5OvVW59lhlAs9
4fplSfaJuJeYDth2htGpMRhgpqJSySWuB49IFXgtpc+/yuXb1JyQn/8XfuL0iQ/AR2E5yqVhtraT
KoKgQRFTmiLNFHe9w6pPgBEz3eXP3Bur4jGJ7kGvauNYAxK2M21mmoA/LXqNCsynguvRwJfDevpW
6xEB7UQozUKHnYnYbig99OI8BkfxbcojQAS9kVmxBa93q7egUgIP37Aj+JNmxzCSb/BZ3TTtuNgC
8QvzL9vtn5IMMD8oq3N7PGuqGQF2FYhAX+uVqWOPooh3YuTcM+JFwTu3Lba7oJy1apI5Nn+TB2If
f44GpLUIyIsyyLbQvF3SHJmvRs2gGy09moFlOsZVx2EFUQMylJwXojge00j1AJZIOSShybSMFrPv
JTkriFutunc/a2Vwm3k4q7zPFzgphBOi5W/+5LSmGOu3A1KsDFY1gd8go1OMzVzE6h61N2d6SRx8
cLDbAp2XRBOsNJ4o0sk0AIdecqvQEEOx5iXGeGjJxjhzlc/iZSjmVF+XzvGNHShsVj1YOy7AA2uH
ownUvWGXs9jZES6h+4eTIsZJ1lI+k+7ouCpH0qCFCIPFKor3F0EwA2hsPzXSKIFw9ykcSCGHdrqP
efH355SkcZavVUEO5O6vv6lN6Xh+Zra5y46+UcMfYRf3jkQT1Nn81TZYi/iW3sINcSyeSpEbkBu3
4c6QSnD/bspebZ9IqvfzSIvbBcVkE3e2K80dPVESAb9SIKfx4R/kfoXHKKKsZlX5d1F4mPde+MoX
AarxdzPQ6xxIVia41J9YXjhXKfuXmOoBkCXNQ/X1kAp0RNcAHPf7EkxuYgcDYx6QZ7+30DJvt1ez
Iflu8iullM0dZEdn1c4hZymsKtpCOVQ7yNALokwItkz7J3zq9oR+AaTJ5sDKkCJJF4SoJ2Cu1sDO
QsycFL+QCiv9nNL1tDe72ZVkov9c/r7iWC2du8+zeoxUL29ZTe13NrII3CcNIVyE6O+RThhomb5c
Ubl5ryoBK0+/RKKrtiQP8ncrXlLst2B8auX7JliuNclaVFEfBtWPnyX206YQWuJSXp+b/NZzAJUG
6Waoox4dQ/FL4LSOVNNY5fA9Gg3Fet4ZfCKEgD4JvYraWar04786dfpQ2ggVpe4HVFMwyLwHTyeM
szPBJ8LieOzn4rFszPME5Obk55NuoOBhq6pcOP8UGBGzpfQM89jazwiGPgTfFum9daYwvs8eCMM1
5jJgi5/UEvodM488rDbMMGZatALKv0qkKs87qAE43hhzHaaBTbtyiKu7U6/8aDBTYwJwf0dgS23W
LqhSP3otzXoJOl7lHaroXNSaVFCmh6nuO8aPrdaU9IkNXJH8q/I9WvhxMnJ/zOtNzxq4OYti9DKT
g1CjVtDAS19Z9+1XxnzlWfsFfCWfm4O1bvzReuhgoYz2RD93lFA7F/VJeDLN6jhRw3Y/nkDN4EXP
nyohR2ZY4ANx0vf1+7Z4G6Ng8HV0nzeQNB5Wf6efrF0kKxBW8E1m6O4eLlo4vfj1X+DcO8aR3C3p
Gblu/y/GEtUKztQpkvHkI6QPbr+EaIgdzgqJwmL0XnfSUnidwnX94vh/5PmarWc/VtNbmFGwnHm0
k22joj4Eghw6alb/gFowr36vuTausq+o4xLE8eiaOO0CPfyc40JmvTbpRFZU0kHepRlsbQ/AvwVT
tD8CW7+9tVfEHuaLJOYBpL5PB5OmPRBL+rw0+GSv1JDVgft+1fed4ZvgxgrcRLo8NmgcKGVnrl+G
w9JRWL39tjQ9LkEdRRa6TuxxRxgxbF/Zqu+RbjEAAfsdQa/PhgkciEGRgrFLXIKFNEqwSb2Pwg7e
+D3ncI+SpIT9rLSmyBSbR9FIWiLDL8/RL9z92vnVMDQneyBnXOstmf7/gr0Yvbi5YWE7uY0hdAjO
q73sHl2xAVk6Iyuni0E6Gognr3P+NTqsbj+S/GTOQhFNtM2E62UYWDI3B+D4LRw6ZOo7hPV/7gob
BOb3BrBqm5Q0q+G/4XMCgsw7pnB8JwwHuHCQm09b8nyuPeEjAUt80fb9VNOAUG3KDY8B9iccTdUA
plCSBFg0SGY8/2G2L+rLRsWVuuL0BMUdtTMHVteieuRKc+tIp3bQAZGPzK+tHXGo4OnEGOtqFK7k
b0MHFt+zSJWGd3fKQp1vPszilmHZKVs7e9wywj5MWcqQjAf4XFQugLluNCnUpKqdwQB5RWEuPsl5
0GhymooYDt4i+EZRjpOk75MbyEBxbUDsGkdCd7n74J0Q9SAwkduXhi+wMMFqaZ1YwBpy60bR/KC/
ARSu28wGfIhsCFDG/Ea52RFU+Dhf84HVwAWiqanxSp4n3bbafMj7RvGRmM9iv+IkQIqOcX2bkxsZ
50vjjRmbmBTVTJI1sy5+n6R1wzM4Y8hV3K88eYhYvzT6JUVkj0gsSdbap4Turblhriyw6yba44Dg
9ai5WGhNEbK/94onMo6cSlbyYwS2PHk1t0rMeP2FUDgjVVP0SecieAcnqPSTnNUQAkwq9/3Jun7u
B/n8M/vbzJv9hvhpZowSHT5dHNQm0G7xe+0Sdv1YUnTUVA8rtau4AvGP3tU8x/5aelOGJXdgQx2p
hrhwRZHjyXfl0uJoihneBxVcPC9NiS1Rs5GwQ35LkrThhFFMgkoafr+t4fVO/v3hZ7pLNeiAV7z8
XfKG/la7L3bS3oXzP0fu7HwcEZmHLd1mm2jPZ999Ohsgzt3lc7zrWD2XO/WmFJsbQIWgVDzQZjbs
Kcuz598EugOIBuDSLRQgeM5vQAqT0PRMJwcsAXJRex6IuKVnFuI+dJbSC+6OkhgJICcgJO72UQJn
EkYWEJ/uyLrCMLWkHMQRslN0+ZkGwnhWfi2mB2RgkZJvbeGC9lu/PVcA9QRCEVkoTMDUtxrZJ0vk
KG2qLgeimLwq8tiNTLrzb+d+oihhgieaLki8iYH7liMqIDaYSMQsaDwmAFr3k4QOGovtEP9qEOxK
8XwFWeUFzuVX+h+nChnESpqQHcKTdXf5vXceAKUhhGdd96YqAsP7fAbz3ryIs1Og7Z2G4JyTZgAT
XVxT3ta4RymwK8xayBsaPFNtR2bVsdmXt0yqxbNHz4Bi5WmlqmumMhRa7n030MYf+sG968XTg6WU
MpAOfwCnizmCzvyms/W60f9ve2kZqyB9RRJL96a4HacdGUjoXsZIv/Gb1x0DC0YD5rCghBmsW877
8zv5PnvHOw76w2/yNJ1QkUrLj+PUun78LhnSR3bedq1N3bQW3OZh5EZqQIQn2hvQC5Ke1WntSy1u
ohLR40Jq/fo8tyRrJG7z36zC/zu+kEdcHg8N0tWkadV8jjPuwcC1Z5ZHwmTNR8Fgr1yM7ED0fCgi
W53b5aZM4fKSiaSVW2jExudFl0e9HbQR6e1w+tOQkQXEeau9kBh2r2VIEN/ZY8TWvyAfSYTIzt/d
jgg93hOJXLDv7H/8EuT0l3/JMoj/ELNbuz7OoZWky5lQsAyyvQLw5oyqQ1qCfYhslCMFKRw1Z1hE
XlJn3SiPljPBLbkxyRWjpnF0s2XsuqUukhqZsybp75o+MS5p09ZeSYXKiLS+2lCy2p31TNdnVi8X
xHwU2szaNhB7EOI8gB5cdAcnJ/x7LvsgEHS5LixkaPNOVOFGDwO6VJJLH/ubrnMvdvzaZTWL8AQ0
4AOppXpNwyJznNNYfsL556uh1PHmk2I1Mymz3CIozMIQol+06bcS7Nc4YxlIBsMbhN4M/PJ16xRo
KkWcTMs9/RTRsxSrEQXElABtvZ8iMAcWK81bZJNbUYWmebkglUBeHVN5DkvTfovPSyWmd83Z2E7w
jdO1Qj4QDl8FrG1eczRndhMh5G9YFzvk2+esXdrRZKp/rutHna8+lrFKqzicsBzzIKaMwB8SVfuj
lZ46MHemv/HJbhrpHEWcFK6qzxYGpndIvU0OSHJWWqvVJpbT9ZEleSHPiWgWLzS/S8Qu2gYhcpvG
m+tTd9pZ11r08xPKUGcUmrFEUS7zgW6mEM5NDt25ZjyPBKW2/SYCLH4/iFlYgvNUgTtW5gbXGJup
TZzeDZGDpd4+NzVOgvmoid72dxNoSUVSC67aMVZZnWxeZXSon4uojodnBnVqnI0xLLcijHIBijJy
drRr/MF2McV9BVfKkCReGLxhRex5jRc/F5zPyEBla3Upg8YlOKqmqc0O3OFNeB9Rz/PUY7l4l6g/
EvS2rnar60iXfoUVVIk5ZTZaAjpF1tD0Ju3VyvoOETob9vKu1z0ErOpu2WeQWUfmAaEzCVm5EAiQ
L/qwJxzYZ8Gu0pdduX3LNrWD+0ky3dmMbvCfD6OZe0IZGJatce6GaGKmam5PJ9MbRoRqhDJioouK
wDeWCQd2EEnxJyfICCpd2XjRl9YFtbIVX5KnofoiFHO6JrGFSqHm9a8VoESvjan3QYfbSftGWLQw
PAfq/Pi7/nEUedRx5hlPeVXUV+CRwIy71qRUIDMcjk+qd1vq4l2KL2uSVzJ+elyeWSwYEsYCntmK
hzR5xHIN42v32A4VqzfMAg5kzr0H/Rm+WMrvuUF5wbVlxni7sBDItkIB/pmiZsEiv+KjLA30sQTA
j+bCa/Y/CnaW4dovQRNlkzRa2oqP/RpMFaONeLQQ2DP2HtVCATQLquZxyd2p8+bsnTc5Z3d0dIis
RgQjKMl/FHsPf7tuU8l02BPOsLNl1mftVc7+xn5yBoleI+4S8UpvC3FLh6pNOzErYbKKWgY9ZOM2
39mmwEZ1oEcuzsfHcITHaiaaYlwhDf76PTFPwX0E6f82X0l9OzXVlEtAX4JOjjXX6h1K71sNKXlt
fn4zaPpwXD4pHcT36P1ffcx2NPRKAxKKLr38g04sw3rWw7DFYEM5QB1eTaUx7RE6uTcMgZbiLTJ/
uZQxEeOdSSYzu4grCvhfnz+VsXiZ278rVvUmhYh0Dr76U9RlkjTzsgqVgRGRAiflXvEvnTRV/jnU
uySkmmxH4mQ3U2AxwkdYpcZ4bIvNm/ckL14d1xFiQrkYBPe0gvi7nEoufTICHQl8gaSsN0ChuKsL
5SuYoJgD3hpXhbKZ/lC9TuJNiZ6Ogi/HiMw/TWTjjIpFFn5pvhdjO2MNPXhQ5PiESNrlQX1IkrAX
fDhMauq3U7mXS1/W4TRNKROtKsK3g26x/17l8UxCvrPX4THitVAGvNP5QskkUOE+sTUNrZRuY+7F
X5UjA55UIh+podZra8h60YlNVpneStD6SzJwtEDUSUxqYFnRpfMbD4KcGZW9NVRKuzrma6Xw30wA
xbV00uZugdUCy1kcvaczkmXUvRB4ehNNtTyXP4jvBhxGheTMoP+nnLxNwRLEhHdgq13ktQWSKP8U
O+z6Agd82h4GTuh0BvCiCxjaRmOAk4hzJOZb/yUKY9+8YUETRPBA/wGJ2UYPYwHhpQoJ/sDFD4+9
fNa4hIxTpEaa/3O3MeYnCBoTIMOpT/PNNCo231+s5/msPCnfwwezHM2Ibt2tZPIBU0nRD0q3k/+I
9lvwDkqx3MM3NdjqlUaoh9g194hh2yrPBYD6uMplhMIoX130byDRj6e5I0Ju3W0zXVaoEiW3ovLC
1T/Vy5hWctNcN8NLNy5oPCNajNEZ/2HM4D+RW0/mFh8aCOOMGm7ausfGk0W6BX9SbBeaNPTX/wdm
aKjTwcgHj8GJFKf2PVScILOADnpbmoxo+wKcgMTnVDCzv1WFFsBzIyhTh+RiVBOsDic53t1xuqsD
vI4G1KBxtwZTqB0ktJ95c0r3wLzxy7dwJ658Qt7QnpZB9SOkNSHFrJ8BYVfP4sFrZZEG+nNUqcoA
6qS1+Aaq7Z5BvdoD8bTGTSYMCseNzQpd5kARlRGZXVOQdq9J9Wz9JcSTNvqoOiG438FDuBjYqL+e
SIWnCfheGMnaDd6p1hEbE9o1gr4ajQVCQDdmq6JhMJ92LQa2vK9zXXYaJcWl5FFsPZG9h/8lLmcB
lXV3WS1FJsegqzy1vseFo+EGSGuFUjv70Ij1DsBk+1rd13YVU8MQCPfGoDjCL6B6BvPi3Y2XnqX7
zCv7KqKIFNx8Mn/TNsJpSseYZlTr3COGTdP/3t/Oz3BjQ4NuGHmGrU4y9yoF2gZrZf7Q37IXM/lo
IY4FFfkM98aDNLr46sYBmf4fBVBmjADguG0YgJ4Wn9dbI1oTXS64n1ycxMP9jOa/pMeodOToAj4n
okFqRFy4neWHMtmIrxFMV4o6yNSBGNzZug08m6WKF6DNQLcCGbXjF9XXpk608drqB6nkmZp9ET+Q
xD5OmHZXRypL2D8cLS8Sgl6QNm1voZqS3bFTGUgnbGg/yjxp1tSQGYWB287YwNmpRQ/wr+n2yrBd
yH7LYjoZ7gXoPaeevh73xidTOpoFyXPjq03l0gFplDd78/J32mEP6oQ7+WK1PgacGv5wm88ywOiV
en3OVByRgbJ862P/SfVrcZXwbVP1aiAb5K8cbuT6VzxGRCAROShh0ixjLttl7pblVgxJPSZ9xHRI
qLE4is02H7m8rUlRK/9k1R7D8l2aq9D9JVSqBrD1YSd2t9nenZxsokBK7L0cLQFgbb+eHSrvNgoe
NyJd2AHk6IiaeD8NOjZGtm1sCLhJvZD5t9B1sxtXCtCND4TnEbgt5gBRlYxc99ABYU4JQPeQdLgV
Qw0XsLGswe9mxgdNLg0jHiivxwlORDm3/CIIOvOM3eaJw2F/qyBFJEB72GuK9SROdJHqBiGwihif
uxl1iBrVbGRKrSPg0to4uLkBT8wCa6XGqSEKrWuivXqhJA8HKRu0xzAYE1PWX+3wuVBuzQQhhfYj
4xrD1KZ3Or6LWSB3MyU9a4pFX5Cah6xtJlBFkxvLF0z1C/YL4fyrG8Oiwnx7jHXGkMSlXUXQLI8S
zrOwf6g7JLZhAlOTlhvXVv2R9heZKH/qyGuQIy2Yp7PXIKeeG0YJFD+VR5MXsvuKhLDlmAxadQ4I
U50/Ncjuz5eLoIfb7F0ETDsb1kQ6THDDgtXgK6lr7NCnW+jG8mV5LRtuzLWh43uow/9ja0LHgbeM
Xjl6aplWG6zAtRBuSFT+bhCqKZEqeHTk0Pflgq2eEyFLjzXG2yhe37DqAmK6ZTv9Rm8h59r0ZXKT
rXk2sVqRARrDlhu0ALQ1VWrM7PNFs2wuESZG7FiJSEnUdlhUhE8ftblUOo4mrW06hBlfXoNvnK+m
A+oqW5e745gKX7/awgCuObdjUJ6JV8ik2YMw3/TaGAsNhvs8fs+xV9pjZ7zkrUX3hQ76zmHzTjEy
xejyouOLzSblVjcN3xmYHMgRJbEYCXX8ozDADoJaivqHjDEZFvGOXt26nSEWttC7DmXTYy74sH3i
zywCu47uPxlToAWHwA40UgFbG7XQSmI1788Lkm8WFbwIvOtl27DpHEs21KzSxazP/JFpkjh6e7dc
imzRbZmdoiT3ZRMdCcCcuVeMA3ZMSYuKmKtPOEfCFUOAcO6YzMpcOMaIjPDzWKwdF2JKzkWkx60t
k/KV0VlzSiAXb+n7kPenUIo0JKpS7JWt4qu1OQY9dcY9n0NROncCb3zm1L3u6dhD11Jg0ZMO2KlE
8C51AV0nYKohaLeVU8uAB/qxKhbVRfTtxxE4oE57nKb7ndOG+2G8DDX2Pr+uNCm2qHJ7ECdIZthb
rO3SkIaSrPsafB+xBwgCLqnsCF2Rfr169RZktt8WPgkhfgbXlt/d1qPrtXm5vHa1WkLJipz3T6qV
jMUX9FHJxrSM506rTmlpzLyoK3j72d39tEh2ALyZoG6Ik+Dn3ZZ0b/r3TFWve7SFVAq2jXlH5ni4
ylTLmEvJm6aD+ohTr6tRfbmBHo+5J4dnuwJIsgy2ka0X7A0eSjteFqpEj0xylNA4zr8A9YdbGfNM
2b/S1H3zVXoBEet0hwLOs5N++yWmPo8I/9StHNqcGuxDplhgGdGwRPDQksQSp6mELwFV0o8p45e2
xgPhlWaNXOC5u1IGZAUDgEcA7M0QcOkLXz/2IuqxJyoa58Z8ARng9DloSsZ/qtwetfRVlMXDNaLA
yFhFE/CcQ1zgjNvkh39E0GutyIISJ2lE+VwkIeOk9B1/jFQxD5IfOgKxu6e/CzNuGyxo6t5fcoJn
L8vk5kCqqIX2VRT2xgeTzgIRtcwz6/y7+8zyZKvMZsnpdMpBXK4sjFS27qWK1vn2pnenNrDOf5d4
G5KT3TKlRgaCGNunBOtxmAsdTQF6dc4z893Zh75BNhmPzq6Amrb7t9umjOnGme1XQORKAtx1+3Zc
YvKkCiq3Z/6/7LBMuOuRKqRrNHsmX5CvZjmq5FmYgBtQgpY8unL5LnbAZjrpJG6MrkjQ9sdZeYrU
iUxtQlLdWO4SZ0dH243YpMW5m1AWSw26I/JsgrYOP/eyK+wz/qdxGgjstHPwyxGpBSSHc/0lyayj
xNMa5v5b4GDyFDSIwsRLYE/eEWulGC3MJDXMU7PZeBLRZN6uRLYIUSbv7F+XXNSw3chpqtAwyPpC
t8K8mE2t/y+LF8sXZS/IOrjiPVw1ZkDJho8Wwy3+36/46cvXXIHABoBiKFdqQMcGowln+wmIrkkp
NFzayA1hpLe6ZDup4GCXIHCOicdKzi6aIMOg4xWqfbZrEORNQBfmdDUw/Z7qwYvMa6Y+H+sKoOo7
+FV+NfvMMzro4ArHM1+DACQRXQKfGDOBMq2QhEH4JTsjVAuaYTmykTW3//qgk9diKzRKSzYkKQFn
K0Abc1g5XS571rTdkqbfE7NqMYSOvzx9Ydro0MFPOcIqGqQUh+FhQYt4/TugvkW2RrvxnXGvJmUw
9CKHQO8ZHfCi+f4z6Zy8hJTA8VN2XVaZifAL9aOGNHbQgztd1wcDejRfYbsFiBQlTLBsBj4CHOT3
RYuCOTTDG0CXOGeFUm7JNzOQF+tQeTl8FlLrSGY4M9AnWYWpilteqyg6PaJqeXo6NCDcysShj9Nm
IJo2o/yPxnnG6YG3u7QSa9sO8CPFBCnDQpy0sYRXu+bvQgZI9KhooGeqr7qBsv1WOsN2P5eZ5riS
70IjjwzczPPtFOUsHkXvPpP884E78OMlxlqU5q6k3HRax/jRm7lKlbpEbx/Q4Sor3tuQa7Y3iFQp
+jT1ZTgfpqlqMd+/t8rgJCEMofV8esMltpWaoEpGGz3CYqp1IlAHEZosN+Nv2W2TtMCzUAF98DSi
JlAtVsTo5J4Tlaixst/kbPQ0gFTrkUJYX5zuLi4Yi7KgUY3M6zyj6r+bwVXsutFFdDvyqoccNrFZ
Y2IgGBzxBd4BxxnKVjfmCxpcxtrAR1KL9LrmEcHd66cX0yNZUHiDaBDddtNsjXthBW/7xC0ANXsy
XGyfYtSTf2u8exyrGbgRq81Ik6P5qorfKUl9zOTl5AetPR94CgR7G7lHnMfGF1Ej49zvbRKol3WG
IeVJCRaL4ilhxBc7LVniiVAQL/W0va3Ips/Km2QBHYu7rrYAuMe+t/CmrPinb0VCvr+oW93Gl4Vo
APnj+u9PyRhu1ndZhgpF5OkxQdTUh3rEv5W5MjdflWs6ooGD9DRbJ1ZHby9wS8Vp8WIx2MIThkDl
dyw8pnI3nnRgXNnH7rRJBvp/ILJ+muGvkngpxjH9ko62Humu0FRqNLPi2FpByWrH1EH5i3WSLbwB
VrLONSnmZp8PDwqU3wf5S1r3EMvesBaGsjB05GxtK1qb13J66Hd7JhqQ8oyff6vLwh5l9oy71/A3
VOl9WxEdNgVHNloyOQ4WJckB3pTQmuJRy0rpZquL+g7jP7lYje7aAOLe9Dupv3cpyd3TJDNkwv1u
SbbFJK9S7wbtLiwo/olBCJI5OTn93bVRhtQMeeT/LtaYzKCC99hqcuhha4M4CE8gzD/p9C8Fhxha
zmj4ouA2m6iEhmfaf6Bhmj+As769R4cxJgteNwKS9XQiIjd4d8xWbVBOsc14A1QA//f8H9q5OsMs
vbLtn7QuivTOpn8IrxNZKKvBg8HNLp/tDx/TuTRsqzbz7knr1wPcQ48P+AZbgad4KKWFZWtJH97L
5/0KC9QEpG45+PXd41VnOiEcuvcLN5gzHbcoRCXskJ+uz+Gf5G5cwt90JpZOTvlb+vt8x3Tdhtid
ALW6S/Fmh3LmltBV9zmN6qtFi7Wq6WTAMgnwRGXUkvV9lzZF7YTBp7u8bgSZg6U/dudinoxu59HI
xSof5MOsA1T3mCblFvhlQMb4ktB79z9R/JyT2UAgiooLlfAQsfCSdfiYC0PMTdTD0VZ2gghJwXKi
vGzkueg+ZBxSfpntY5jPUp8R/t0pqZq0sulFh/sPypEI1lHHClCov8SdiggppwA79vFdMfSSJBwj
oGMhxSXVCBsOR2RRRQG4yNLPdPVmlWoSsaBslLZ553ouSkxocHUIDySPOT67FMfrxrtxMYFHYpaH
Xy0ByUmg8M8ZCFRKThiGU+BNJvdlSamK6iUIWm60HCdyawCCPTVA+9ET/Ry87oJx+zknGKZMVlhk
Am7H1gYV5UkvpZ5wB0m3vfHmtmMs0JYGaQ8YZbNN2hhyoojT5D+Y7xL7ha8+/6Oaa8sN0JJOpHb2
MvyqfhyoMNnuOJ7P3IOcxpVLYJTrbue66vkS+oy8dW7FiJb9bKf3fYNzN46OlUe0b98/RGAfx+Up
4SDf+vCmhzbboQBpgd1ZHHUNHz6q8uIHHb7pPCeRRDqmGVBrkthAxdWug40hti56ezqdNzU7H2gs
ACpxHfEPtr70+/JgNzqAY36qAML9Y1h3pVkIHavlEk65Zg95TZvI2/b4YmUuAqBJb/lhd118IFJQ
oWgTkf3kfCD+V5pEbhhmyG7R6cu7uxz6hg7ygmaLYGoe+YVYnrrj5jneCEAbb63L7E0GAjz/10RE
sDS8tvfUvPwtetUy9OqYxSNMsz6Lc77aUFmHAjs/qbytg228cF3m8CRht0+zYgFCndf00zMrxwRf
wdZlJj8lUWFeSYWV6NiSlJK4S9Ir0BoDISmQCgMkfttIutt3JgLtr7ITywIryCNUkEomW9fVU4U4
Ly+Lt8CtiZL2pcK+ksRx4foTatdHqTOek2MbWo6caQ9Sq+2+KJOF+n2E9tk4dUyc8T9XOFzJr+qm
oYVGF5alhdTsiWX9p5Ht07/FZsfe4eCGrD1mGm3o+6Ft46BwdkxW4fFqrMf/d0zlLm4bd6eHSfvO
9tzPFUvCexzoiV5+nP+5WuX+4Wk3p5+S5jZ4r+HtKi1oFPS2rYol+DjGCNwzhUOzDaqLo0vzdffJ
WYjXQyUlwAa260VKeMJWcoYca+3GYdaDCUeTyt4kwPpGHfuXfpqOIiU8VcKrvJdik3ET+SRVB0Cu
wLqL7zVB/G3MOfQcQXPL6Bj0DiZOcfrS7QzQ3Xqt8F1nVC4RTljD42EjWDwSV5ukknubmslTLJR5
YnUXEbSfmVX1f5X2SqIq7VvnKsztpTISfCve3H6hFYtANk9L7SK85DJCF4DPij5IRh7D9RtHu75V
OzPArPIOEcLSnAnS1VKfiZ6j2peJdjJMoZC7zPdB6w5Jj6SxnpZDEpYhn6mEfYCKwsq1DcdmDpBI
V/REmG/FYzMTn7cr1S2yzrYLlOoZDCkNR351TJIbxatamPzYxSR6MxLN2J2PmUlUaE8nxxwKCBtb
E6e76p4+wCBWgOH6y5w+2nOZ4rkaeMQr0F1uSUN+0yVe5U/ccblDugFTgTfNoooZaMZpmkAcREqc
8KCBSBPsDyP8ZY9bOpkPwozk9hazYqFYs7MPCJlhj6XblJpemabXTVXWtSWC/XFrfKU1ybSUpzD1
LmgR9hWlnxKK1CVOaBnZv1qFfoX2PhvsmhWlgJjISztZbHBGpt9pyTv1xPY56ZCDhim343GvfSVA
osTrv6BzLovB1RPk5wik7xNQppJhPPJHYl2eoKlYquenwJ+QmktJD54M9DmWPYCwMhBm7pgmjXSs
21HuXhOLAWri0MZVhDy3EQa0lR9lesrw9j8VzqwicKkZu8rXMmis/VbylQstpfWDQDRDm/Qtoplc
s+mNYpBg4o0yKffKtsRtEfZfIiReeJxVdM5DTX+ArGgx1sh7KwR0SlNbe8zFvCrRPEcRrHRJcUGk
5adEhY7Hz0QbVzPNmAyWN7WhUjx83W5NoBGMjhDQR03N5cLvoLqGHCWgjp/OD/CuPdavQ3jBcFJC
lqwCG5LA4EKcFVtofnLSU3WDeNFE5bgynt3KfZ5Z7nPt3PGIz4+MGTF7JeePzYwv20Ikl90ZFgDy
fv7ZTLHoX7w7288a2vf6QUDWmaLGAPouu8dL/bBAN/zTUACbJNWK7BF4oiOBfppab3T3ax4cjUEa
pehI0zWueq8/g6qQdR80oN2P5fvPIpQFD3iuCBbCPT1v0MJAbkVd2tOVOz0rashC1E8ZJzJIy+Mc
rrtEX9RPunh7vDBYud8FdIBn1FNyX71hkv0s7uAc+auDaX5ZuoAMA35j88PLsyn4WXXIHUUJQxmG
l7FoDHMONHW40WM+741e0UaxExZG9j4fqIWQhbwaUCd4eMRCT4SdfVCf7HykHD5vJRPnmLUMh6F8
rxnXHbteiHDx40yMCeT3iE7vK1VOZvByj+1fDNM89uOUE6l5AIQ4SjlS4971U60plzu/0nB2/RGt
vUQQHwJlre2f3XaWQMJTW2yQpobdBcKRWo9lclCaK9jzfa4JgeL8YKAEIxs5Vhevjl5vqRXUnNBj
GH/AMuBS9ciHfRs9miwhBxJT+didF72QQzzxVRC+cGB+KL5LzFWPJ4uQNE4sWb/3d0Hv9lAJuy+W
LbdNcwW3769rAOmdewzkBTwSsWfGLWs1QDsIrT3fPPO7TI29XqKSStUJgujtquWZdZDxqe6h1TQK
c4/cl6aOSpTYmgA7KrBk9bLQpC8b8e2amepvXlZdqm8g2KYPBAMhCpir+k/+JNGu7/6/b+F7YW8W
5PL+/HhqyJMx6fKEvd3FkW8LJQ5D2889rGyAvf6ef+igFyDSKkoQQhpD/SYL2bDfsK7tuuoqu+6g
63WM/f/Mrl+HyduKzSwESr6fdWrDZdQ1exUNbO5Uowy4ZhG0MraOqnNXTKWGToP9rIScdZc5w1Fs
M0Y6zbcL0duDrl9U9/Nv1WCDJiLxGdNcnBVgvOsywln72zshdz42gH9SiSL354HcyDc+muRP4FXK
imuZ5AcPxEToPkQjmt/8C8qKLdWuHbLKfAqnA55zblmFWtXRuGB43F4uaJXiW4cNZ63BjVrDsyOH
dwD0ctFkFL+DT39F/JB3PSgXc8zk1IlsILR056ZPKWEsZF0ktQw2pB0TIx5jCbCoL7gvaBwCN4r8
V6BQhW9CjD+4fWop220s3tJ2zReS1T4WzzU9BfnvdZeZ/qrdbm4i1lyLNQRlW5Z3MZ8g8qJLodM1
QpCy/zzF2v+GLpuzVnKDfChmwKsHzHoR8n/UcvsLmSXvYgZW+TFsV7w8n7/CH0jF+nftjMcfO7VO
pEaQeV+tROSDry+7pWXZO2kM3wohAJ1jJa8AcGNhSnboMLC7Fez3gZVvhiqrJeljbWthfVuzGqYN
lEgZ7F1GvwBAkK/M3uXdPmBGkPnqUc4Zy7OsMBbmV4E9/LmiyVfoZMcuzRjK7G6KjE0RIfO586/h
SH5QRrr96B04SrdhR6L9a1GE5/xNIWlr6uOh2WBLhZuvFZAl0K+hBUaAUbf8ZoD0xJJuNHZ7IcZw
3yM0Cp/t1/pxqO9rta/qc09L7A3Z3YuXWgb0d9Jv4Ykg0cOWxMK83hEupTuX/BM3aeUUa0rqiMHm
a0y4JIr2hOPQY34uA5IIbrxPWNl1qf7lrRRulv1NYeWGFQhnLcDlJvMHPWWXg8FregkeXNEU1Q07
WoYx/xKOrSamn0CsgkMxbXNZygw11aQhnVGlhEVyXmTZnoDckQT4zrlEZGJOUAuxgl+0QdpbDvwF
EDHs0Q9dJ7mPrxvjmufPXf1qpWAzVTNMD6mExctuE5bU8SnPYPsJ760/EYqL5rebESOZ1fKCKlKR
EDa6adIz0be1bhlV6zhzviCx6A9CfZcDsq99QIjFGorqPliluDl9y0qX7p3w2Y/sybvp5+fpzoY3
4K0REKNLFzs5KTXhlxbrJ4C+tAYOFGtIkzVerKdR7tICKqAap3fBqfGk7VaB7zWRta/rzgIEQVUi
kHrWOpHC4n6xZtw7Ypwqxucaq0IPv/13EgIs131OSBVKv2JDMjoXw4uQY5UYrDuXXfgLaXOG9rz5
BIT0Vp2E4wS6BgaB/Rvd+FabUzPMV4u0Z7ce59IAzx2G7nIagq8iaZa8pt8zyeVWTi0pf+2R/i2b
uT5vOpeXBZ5H6zvW9FG5hBV8sNSSOS+k9PcmcURP5BuWR7Zc4HsxGJh3Wl6vUxMZBb4LoC5Ckyxp
srTAPbam3FybiSRyhk3W/Q2ty2C7u4IEm3IX/pkehcJ3dQ5EcQl7e1B3/0TgmljTGr1UN7zU4fHC
xR8POTiSvV5R4BjCIREzDqusUAlmOWfB4I+88QUjxima/SNkdmwQlSqQ0A+2Hvj+Kk5REXlhXI4J
SLSA6YNRYTOUShLj3ehoHOxnk1+o9uGq1jP6hQ5F47nMgPS2NDgGzDo2Zq6OHwql4MoZ7FxIKJzn
rfm5VquobdRLQBddqVFPQLjCfS/PBL4cbdI1U2qWxhHbHK015HgeUY45Zw8Cf28F4ZvRERGTUTR9
eyyfL83LFMEg8CYUjtPSSyaDisJLpe2HJDqcMbx8YU05jUax7Fe7NZ6E2ADODIPNP+KtNLEOXoKo
o6kvMNBAhiG09dzVt+agEDKCrtPWypzQcFKhCPMsK0IdjlLSkYjM3dR2tjr01w1OFBQ8ZeDb7Tlc
AgdHWAd7kZeaHPkNTiKkboh8HnOS/TCI1TmZ6Y7KoFNGrv2FI9TbkMWnqFuTgwyLSZnjZkUPhRym
EJaz2CkoKMAG4p9jHUrZigM5Fe8ggfofqDuIkjAUAMD5wVvfVNIJv8JbR855+H5kvXuK0NwHBCTM
IvaJcFLil7Ez4sA4O7RiMgySsyHP4hWh2LScuDCkGD9pBSAwJhWF8E9WQSIe3O5+II1u/ngCpAtV
Rad7iPnN8guHq8kc3ikv3cXp9gCtjQy2Xl3en9xbI6Eniz02QSFjgGFVy9ynlPvICljQOPCY4C8x
6kqaj8Q73eEQBmqwwb02GjgMQP09YjGiw9UVHLqSOZrswe6v9YdumJ8hzCedx7CkDN4LRqFfIhzB
kcL432qKIgmW4aHnBKrtj7fIS5H1c8QFYboIZNM+tCPcOZtVeDtw0CORJp32D3VEK8+Pjtrb5u8W
+S7v19+x0vv1jI2GoxW1TkZ0iqRiYWCfY5twVO/sLM9F50pedPfEZXyl+U6ZO6q2SZZ65aC4zf6g
dQNfhmkmGd6c4XUzR8lcf0N3igynAFxzWCGVaKhdQHGUT19+PPCEzwU9Lw4nmTkC1ldewSrA6C4X
mPHccWJ5aoi+6P7O8tu8IrI2/8ZYSSG+jCOKpdo18QhneBCS/ETnbfRbm3fCg/nXO64wgA7fSypE
dtVXgYBzPAFke3MmO81VWCxYqllGKYNmL4N+YHB8ucEsTioniebA6ZO0cac39ENessQJo4cjVRT8
8PtQF7uG8wk8KmZ9lKI4eXzvDhNrXlbrNyW3KXyXGufNJiFleBaYOMSwRjRWWkaUun6CVRFO9qsM
vR6ZRSZ7XDnpvhiWpNnV0WjtVIJ/E1GeH1oiMgnyRUWQRk490ayvPzUkb1PWt7kVFcC2dSIK9+kh
TCMCoErxg9Cux/Kj/8p362S2gtUlMEgsOMuij+EVEO8d+sVS77dPYWCF3tZ12MFOuCXtZZ+fCUH1
01UgYgub+21gqQ2P6UMvS3AuWLLMcgpU7Ympc9cOC2yspcCEwSEtSy7wzz8UIJxfdSYpwXzT4uVJ
TugkV+jvgGh484eO4LKzTbY/jKvre1+moVXPzWev9Y6TyRlMwkRWKnXh5bFFYb+sECaiaTmQ1/CS
EAyyWC2G+zMqq3PyhJmt5aFVxVFx+UFF0/dXG342NQZOPF76saQ5vhIZtVQNW7vqDPvjBJcypjIN
UsA0Sid2M0G4+vD3WEddgHx4ZiEnZndYfL8gSMgK0UFB6dBGVn1qftVEsdg2PGmgyhsF9pU+9Ijz
xSS57msQ4QZoYKkjqrH7UXGSsu06N1iC4iAuMSsP2g4cOgEOWw+BARbBeR/6hUeuHh9FhZzNgXl5
diNuVby9z2gkF2fO4HJSehbWdGOez4MfMVfxU7eWqtWgmE+HHnbZeN6ChCkpUzeg182D16mjh8zF
CxQN9tTtmcg0jRBfnSwN97/iLQ1rhl7r09/bXJDXc8OP99A76wOOCiZO9KBMEWFqvkCCJM3w/R+j
hFM9fc04ngPhls1fFbFuUp9Pj6C1wSgSNIDeSYswD/fMBAoRBZPbXbfmPfDu9t8ARkXzPTCyaG07
KN8QSSMgdH3ZXaVPVS4xK+ySAI7u9sAmtzXm7/H3BMViP95dEo26njSgQBkD/XtmnRXXDz7B4WK5
HKTphjDL1Pqr/yxp1yonCy5AMgAJZm7FQXuzSARFtO446YXhoUUtBnOOjoGmEuXrltEF0aIH1T5y
FFzBUj0MYgZsyzosm8A/Ooqk+CsESzCl2YlfK8pkx9wIEkH7jeIcFyMM9336Qp637zeO5lKOOldH
apPSG/vU8+Wwn0NVPjonKutzWrFlR+K+IdfmqLepVUJCA5FOfVuC9RMExwGdEmxpLx8ZGisduAe4
UGMNFXnIfcMn3elJtvm137n+zUCQ0sEkOy0fQModYbhQaeQq9Gfbw3V8sGMiWyHoXtnfZroAkJbP
NhI5jM1nc7HPBOsMCnTFe5QK6/uUE/COyoBTyArOsB+sQBNbnD13XhwcjU13m0F8h5bjvAf9Bubc
WOGEcMWnAjFz1uA/zEv5GfsqcJOJAJnCPG/sGErrwtulI90y4Eef3nZ64jhmtn+x8UL0AfwU1fb8
3VmdemG53oP1OqtGBsPoNm9hBKOoJOuHZhX5PC4sPTNcJ3+654z1qx4mufwKZ8HchjqFVB/Xp3fW
18VUNil8YAH46F0Es6DuaRY5i2n5wLVWeg1b2CcpWwBKxFvoO9XK355IjPOkdOH7gx5y957KZDhP
ppWfTXER7BvHgQOnFwsonXqpaHu9DLQXUTlrX7S2NBlsgjQzifBbZDX6p2zeZW3LBYnMW7fUbBwC
xdKoK3/Ti0BHJkwHCpNNhyJN4JzFFG31ZJlPsa9jCeBBVIIBtDTzLQYcsBhy4xTeC6iGkwW78zPm
q9wjhvBCFFsrCVdlf+Zv2bzuDDBUqDHyXYK3VbO6foqNJTyeu6nKTqxHVxNt73JzUZdBcWmD3yIO
ewlptMfmX+bna81mt0C1+JL1+PRnLsg4TH7fHFcaM1jo1j6XqiNv/gmQ+RqY/dFcT9z7Ds48VR/1
BUYea2/HpsKOeloLSA0mSbjYJ8b3wbXiYxzCXluXf9AUh9guMoTrUJ7PwQXjTaBGgoyZR7LYlG+V
Pv9BlveK7TLgVneCILYmBe9T+NtwsgAn31qsC3hIJSkxXzT3TEsKJ+JOTYs3cuOm8ugE4z/1WvZm
5CR0LFmLYaeENJhU7WlhsUpatC/xeSot+8LMUWkFgHVrOF5TnH+uSgDA5VXZy8PzFi61svv3Rmmv
08xe+tea32kmyztYHMEr+gDh48v3KZQANOFoQBvb3n3qC4Qhw36TojjJGxdnggHkiGYWNv3FGkS7
1I1DAR5Pr1Io/6g0xs/c6No91DHY3M8F4v3O3kMlbpikBNzx4tf0oL+LxHU8a5OoW2KxRtAYsR5+
Iex/oToxAuRPgDigY0oSGd4R4Wi0GDpFpViDLlQ4FQgMygK/Ecke7Q52SJ3OFRaevo2u+I90LlsI
jGweXkD8OtR1kEqU6EUlqglCUxVs2zNoUSJnSWmflPh9cFdTb+e4JeuXbFpoUfUxWfPE14PDpXZl
K6qcMhsXgVpcLvOunAp7uUDkz8DRTQybxyM2L9I6ZiDgiBH7PtpLUo/aMFTeSl+1zLflCfBgGbC5
GRBYD7N2O9xu8dgBBy0Nv+m+K29RkTdvwcsLxEgxaOdEO+CXTdYZ0smSmVllNEfLswnaY9q8Poty
teIHz20UfIKDZhb0dOnZZp9AhrhcKyK0guhOk+N8yoizWMsatrGbGiBsOWrxPvy/6V1CGHJ2NQK+
4qdzqGHmkm2uCUWZqjpRgxNtSiXtmmZcAV3BFPPCqcKB9NmFu79BJfPB3ciik/LmNFOuV9HhhFhc
Sd10vYlL/6YO0xWAZo0ICtkAqCsUGTfeWPL8roMXJufkijgfqV2Bn+6zj0etNXno5xEK6NdAN2vE
UXG36v+txZIcOnMFT+m9yx+Fy5E7Wcdy0gCCcKgn8NkzQ4OuhAsg30tV2soJc4ceo5LESQ3VwRL3
9adajuLE75D0ZRg23jUvLb08BRU5JZDnBm6ZFZIY3xgTBKE2CLpvtkKpoSfjjr0yqNxE30ggWKb5
V/3cuBSPnNyz2of9RZ6abpCH2mHYZXegfX65g9M5Ii9eChVmSGodbZZrVP2mgupsYpZ5XzTnXAZp
F8csoCtuo/R8sNUXrKPaQPgfroDwIikk++YTxyYQbO4Tzofn6bIPRvwSRF5zIbSg08NP1zRQWHtl
ebspxYzcCdtKt719aoLdrQh+tixe6I4bSldA4XgDp5/bYewi32VHA+TotVJzTQmM9ak5TtXWM/Mz
h7q9PuoNgAhiUhI+sjsuL/aDVSpU6L3RGeYzzoTziYiUL2P7JTy38N1xPy/2zKhRMisC2ItnbiAW
IsAEnlzPSUwy7VxtkRgVb55kKYJ6+1kO+fv22fYL92T+q0Rq4gSGGlX6+z4lKN/41Pb/bVfDOeJ0
eqAHGUvoENrfXbafiv9Mfh5qa2r9Nft7oDhy9y5rAY+0q8HkC1+VxKvOOZG+3NQ3v4IbjQpVBXU4
jEcQJ10x85H2SSn81ut2fjt8IIgKcI1fGkxviyPhmTYWLacAhzflAzo2KaIkPU1WmYLTKmdV4HQt
JoUmHSGp48OWqJ0OcUejiPjxapoNMLZAJVSDrtm3+/ZbiMMtszEsRHHm7PgVQytv/AY9yagAlhdy
RHzfVhjMzb6ZKDP9sf0ORihQts+BXiatCY4MyFjavhDKM3gHGIggYjNB1oXIszQAdjZBQvetDRtZ
MIBkiAdWFq6SyPrxjnjSYWmWn960PnQzaR5y+6DPDA4m+l5nBdBPjEUK9e8Hflf1UEnvAj57vm/A
eP1F8TiIYDSJVqhulmL5e86pQ7A3SZ6D5Dmmp8s43sWgMS3/p/OVxTbC3UHgX/Wf+3aR041+BbVm
0LtYoPU4HJMuxkszWDycm7F8VodUh+dzhDfveRvwQPNxgdL3ALc/DP2bwv7VA5vhEGDLsHicZpPm
G7/cBVmIdM+uuqaQBHXNwgt9gvUT3UVCyVekle1iJLRNkzq6g5suRsDmKntR4BG4UDQru14c1ukU
7Skyr1XKHhLg3bS2a0ut0KMs3Xn4abQfBQAvj4meW1pW/PuQZGpAUXzXGZUnuN6QJNAErJfsAaF0
YObQzul11ygvHdGA6xLfH0I3izx+jQSOIbtqB18oTvgHzgnj4GHbJpFzOyNALcs74gUbZ2PmbkJw
jBTwHngCtB0Ke9PIetx1kTFON4vjWHAMzfprL+V2cRt2twOq5dtHMS78PmzVKDZ3fkeB0iAPgRok
3t7MIVF4uwk7VXS+F1w2QM3gEImk+bOuYGuEW6Wer5Ga0XL8QNgXeSf/w7DQyGczyeMjfrjrJKiQ
nciVktNURRsFCZLCZBvwYr4f6QjS+M4tys+0TSEOYh8KtBs19+gJSLt4vte5cAYwN+b6VrigMQCm
JTyOgIcJCjonsTcWhMMn+PQskJAoZ6m6zxVxP+KajIrM7lIla72z68CzVrQ/P8Vw5yxNnwE8GX4x
7ssYXbQijh8fQcUlGV8OakVICKFLZxhUS5ZGUEwt1RXgIA3CAfyWjTPdFpgkkITkcl/4+fNpiada
Ds3xgJ0pKDzEHWjlP+3jkeqxbKOt0VrPv961H8ai6hAxBpZmUzcVvW77BOGEQDCSSrBJYNBTSGH0
fxihN3LW8D8vGrWoBzbSo27ObngalxOcvn8Kd15oksYjLuYiAA18gw4drWfmN0drpdROCpA5Mujg
1m/BGeWl6dbAADorwJyLFWOM34ClYCAw6pRFQ0dABX/afbW+19OgZTvDgkjVAXGV3HtmbQIt9eBd
ySS81udqVdx+bcPfxcDR6bn2dTO1YZoDqpu4jbOVSgMMXvJNzHqYEpM+Eg7JEiercO7Xop765nCh
jXwigtxM02o9QmdSDMCIUZROO3NJVjhA/CkbFUk6BJ+JcryNFW29JQxp2ymmIIpEUvJTPs37nQdn
zkHCW4D4tO/1S0zPnTj83ecqw90oXApM2vpZI9B5QUXQS9P9+u0u7fmE0A8RHBPQYB0qokto54bq
HTbrv40slsO9qDs0oiutOa9uI1vGl535ApUbjr+5aL3mqjy+6M5OKPA+Mp3t2YsASTVLFt2P23SC
aGyHR/oxgGP0JSVYnkaQe11qyyUrD4lzQlwNAcF69t+Jy22P2Q4j8QGH3lhejzzzTdmUE1DWkjuG
YMe+eQire348ltRJai31OlwX+Q2WwN4syI+vx2xPl4yY4LyteVZRJg5HYTWm+bO9DdkQ2T5zay3X
NiZuOiixDaBkZj5IAQ/4vH0a5RRWVW9h+DyJLdeHdz30D3X3AU+TP/rd/GYbcsag5PhK+5DUsYrb
w87WFQ1McEz6LgxlOpK1NDvqNKRKZDDUw0KaEfr0CmdglRv+jkGBew+2p5kEZFaPtMncMn0qA3pe
ToIqPTqg850LLVIXT6F9zKZ7C7q6pfWYi7+OWKBHgS46bqXYuvGsCkOxGOYFb3HmNaG5p3F9M5P7
PW3Z4dF0ZAT1FBwRWTsopzS2EeTBPnTXkiQheUsYZ0smSzeIxqJPfhgTXxmMzV4axAbsYLcOVh32
VY6cuzosaC9JmsOB11ZPvT2aJD52TSjmK9cAEty6AVF4zNtRNgnx/9ZvyU5i2Qlc4vxaAj+U0u+B
ufI97tZ/wEfcWxUwmXZB5BwQAHLP28ao7V5N4ILrdkUK2sF66lc8GuRKhnFZRDerlPiyYWXFGk4o
OfTIANgF7+NfLG8RPcJPz8LJA2WaTO52+Z9iPpMi57diOpzHYEPiOeEzsUHuWOHWxDCP9/h/oxjp
bNO1j/aG2ZBvXNkKb32UhCNJLYkPAc68cl+galrTHSXOwVDKAa4TCqsCxoI5m9aaMN9yNBt6BGvk
5CZwfTjVy/8vAgOpLlufGoRsuK+nY/ANxV8C68bEpi4iZNr0izShzKjZPKGd0ixorBSF868c0cxS
zKE65ebDTpGAM14jU1ahGT+TSyW10ipZk3IJ55m/ia/6sLys5RSPSt4i4yciireubNQleRA4fjcM
OmGjvgPOMeSUKG9ypqsfeRTMgNnabInOyEn2KFedFxBUHEW3ien55cJKHYZnCLFtpfZ+7gUqIpxT
HD3uJEQxDTWt4+JE6/xjI8uIySGmfbRF4+v3BJjXBE67QgfUopbPI2bX+sGt51X4XKpW2KKu1kW5
SJ1dz820ibs2gtU4yEMFDpKpzniA8Nw0GAxgJyzAx513bRUtmlhLVmtqLrwNmafcOb1ZoS8/wNeu
FNLGPQfyMvYFAdQJtFkmzP7GxQzHfbX9/DFn7WB2ODLHIq/GCB6iIPHNSldP3/UpGAJ4fwMdRB45
gBZQWG4Y7G/h6QmH9FvVNel7S0FAycIM5qrl7hKw8COtyWBzXWCDNMCpbdnCdGYJrGA7jbWBNAda
SyxC+z3bQ0gIcjnjH6FHSEtbZhK5i6rZvnlWTgWPO30vdLz5OUPQ0YJhFJZO9t1M591NTjRRoyuB
9u+d7UsJ4XwDQh0X2M5RquJ3DxbjMZ3/HE2bKt3b6zbI6FFfB1AFVrBUChriiUvHLjODIlTJ8bKh
9T95O2ipv9os/l37Qmo8LVLHh8cRu2BU0otavsTpNxfChRGB5ZGh60xw8wLClMe0/Gt3e/WOmDoZ
/X8jAKtuuWUXfErEiDM8qZ3uHa5f5Hn28RJncg/7BJuUbsPsh9vh373vyrht+fwBxBgVxg0bY13B
sgGwHGHzVwPqwpCkeSYUzV4Y28HnbWJxboZW5KWmh6QP2ZBHGMkLMZhCSglq0HFIYVldb5XzD+If
8gXWVTqfcHlwX2f1Z+D5DGhBaPCoaoc1IskDWMRfOwMd8Is88RneZcS2hIdakACMADg9aC8bBBE9
V6729jpDKOomVZIc52IHskrnZ8fdcK2de9r2GXxMPOwq6Q2RLMiVjWJWzkwk0RxwmOrG5HOoqmWs
VTi/8dtS8mIRP7mD6ui8/q3Z1726D7S5zxL0rTvtcmYEdNMDTL5HTdTCIZG8DRf3ukUsDt8txY2I
WCf5OstzIxPrfwXInivDaniMMwvCn6ZfOLlNLw0FSrqMt07SKVAbtR1N2QaA0wzc/qr8+ymhp+56
Z8xRQcd2CsVpBo8yORVJMn/jr+agt/+TCrjSBt50/wxIgzJ8j1KXrxSqDGf6HOAKJ9PRHIAIyk48
gztdhJ5pgbVfmK4KVuYGZVheEtemObloyMYXu0h6wI7S+4qhUt1vGWHJSK0xR3YpjvjIwD7o6C4w
8Uc+dK93N5us8Ti9K6mDuOq6/zgCjsT0GyDe33V3KE3mn4zRa1RyWlpkObS2olfXtXp+BV8I2PDx
IlOGE9KoLjOLxYhYnib9JNDodPmhs4SPtr8WlQkhca0TLB5qFvvjzPpGY/PQAQgIrcb9GXRsxMSe
mHq0yHer0P50O7zkFMBWASKcfiOqZM/z5pTI/t/MmWThpFV3Yaps50haaBj0pKc9aVIFzHAsaUr8
bCSPT+mJP/ylXTXE/8UM1RS242HgaZ3y2YSduK4TMY54VcQ7PyF5LFr7kWEBhEmrKwKeVdvJuT6v
jZH++SRhGkPe1UtMQDj5tO0ouF6d20fcCNu/VGQ9Uqkpta2vF7bla8Gdqhmx3bzmWZq9ae0Q9njF
7M0Bza3x/0AdCaXaFo8WqlZ8tqVQNm9moeYojx932GnAQFIt7NVVuh234d9nikGRqFocYWlbQwNB
xvjIjNKnpSsIYHKontT5cSDilc3hFoTalgXuufkl+Oz8I14pwxzeu+AhEgBGVeGrQOzSz8vwgV81
fUES79uUJJ8N5wR+MwLsjKHsNoz8/sz2A4suvGpo/oIG0qdMCY8S+9u50RJbelYAJHYgksIfl40O
k7sbuhviS74ywqBfIE5NHFQDg2g1V9nZ7436i2xnroYStCGRM3gZMbbkHayzK5QqnRk5CJ41MUgJ
N2LFZ25ym249EhFYDxMDr/32gG5tfnxJZmHGAb+B+Hy9O8xWUX+uud8MIevxDHa3Ka8UAuTn2syg
jBRyrupoD6VZ0d8+2rRAwrimYodlPkpcCFYrh12mBera06XaJSoIqd5P/nsJP8vWe+lq7f/oJJU5
DS7y+5MYaunjyj8LKpf+0qXHlKDai4okhPDoONu88quERkM/o+4ZU5SUQVdc1Kj3mtHs4rzJalxw
94Kgw+gvSdvvFQZH1XYFp7LV2S2AdH+lj+Pe6CKtR+NvvKP1TuBN20odcCj4z/wqsvkBBJgDCTY7
Cca5Ep+5cuViVsJtaVXt/iIppHcyKFs1ZNrjg69wkW29rBxHNfLcWJG+WsMQIKtM/3f7alaD0ibn
yJEcnRJIJflbdzymHXmoadHGbTA2f4l0cxvmAwiw21IrFkPBSYxl2dL48eEjm33KYTHvkw/Hx80r
a7TXmIpPP9KIBAlpkDIvSyScSdo9yVcn9s3bP00rADAN4cWbTrJ3cItIO4E36/c/wNYvJZq+kw0r
8kgKn82orzRR2+bHGY0Erz1Gs53iuM4wWMMQ1m8mL/LxLTwcZ56W+Hd6A5acoVobmlX1zkpYCVyU
9k6anIP/nVCwyEJW24wl4nYaDLtN74+ea2Wszdzip/aJfexxkzs3ima06hqGt9Qb+469DfX6T5Fg
BbmCIRSSPNN0fxwF6y4CFKDqDodI906xOq2j2WkZNt4o1GjKnx7sZ5ycHqZ38InUl6Lb1+p74hNU
dV92bdSNL7w3hH8oMnGvnNS8NyIUZy/jD3Im9FZbiEXaKnWf7kZiUbSJdLAAKBlaX5uMW6FDm486
DxuqhyjEtkHOzR6J5jUp4YQLFwxdjWFHfsgW25moCwpBymScc+pDHPcQRBKMkfrDahzp5ahK17u1
5sRiJOXnc6jHw9cU9DpML/YJ68g9O6x5BiUdvq1Z0aM/xLSc7y6pnk81G1FHxLSIWc6wkUWUtBzr
d+b5oxA+04OVSpmUkKV63XjyF9dpvaBsFUTUf2oORJJJ+OXX96/EulpNaUEC5vIr4ddMQONXliSI
YzFwDHHkuNqxM/W9fNZf2ulI8uejN5N/qP8cVPmArx8mwM1D1uu9KfpnZPjdVPc9+rQFpF3NjGdw
JRz1S/loI2VWxVG3ZTxGAYBTdbvEQEUJn4TrnKXwND+4teTRGB1lj60pTuOjvEM+QM5iTXOilXhX
X+oCuPsEr/DEX28WE6v4K5j/2amxrIQ60B0dg+pS75cB4eulTSkcZbJgv7fOvxQjDtsIz3PKGTR2
zUhdvugom3NzDad6BmvYIENjUz5j8slVjuKzEzyyKn7oFo1YyfPgpVOilPP6guUsf3yd38ftMSzh
KnNdzDxEbazRdEKCDXL5Fixodqgq2NrqIvCHgY5/KlPRkykTIAIvBn34oCzrykJ7zx7SwOegrFqj
gQaR2LegkniR+++eansCuG0o2Xx1WONxEzuYnhlYu2Z2DpnqExcQyqlZiXQ4PtOS0ZnT/+dBNsDA
9nZZwkd4PvTt4Moojji6KffjR/o1iNu/Z2mKzXIsW5TZ26fLEk6DcGnvPsvTsXgfhyLiABtu40Yt
kqszAIJO+mv3p/hJ912/bDww+NYUf6SttzsDVoR8qRCjKC2gQV86Z5ipywhwDkbQ73p7Z9RzWAnM
NbVcj3YRGQP0QN/q0ry45f1LwXRJVujwCGT4ObLTTFN179F4V77LRd+Agpj782oVYEyWu2TtV2pT
PXsW3ckHWYn6x41fcf69JoCmkS9p+N5FzTnibMPC1Wrm5MkdgE2tLWgw6o5hFlCNm8+ae3gFT5+i
0bAijQLtIuPWRO/hfeWxkORxA5KaTW+3coPdI1/Gn2PisdVB6cOuWxCpk+68stlCCYlMszC7C1g2
cwz7f16PH0QGBVRqjvAF/oEO4Q1pJiwEKn4z2MTUpGmXPIzjqFMbnNJbirP6pTom2ayWa5/klBIu
FhO6mRSyZ9KFsjj4LysX2lFPYLJUjuxHZbycYtsNAYxehR4u4ow91DmDWAMWmGOH4MI5JHzYZKaf
q4Yraz2itZj5BrQX+SYtw/uHFpw6vAFXjNCSN0P6L7f3EQJyQogtXmHY3kPaIIsGTyv5JyH6CZP2
jOiiBBKCiUHGfp4gNwHzTLAvbwPPIuYavR+7mfbnZwyqqCD7E4GSaMlrduaHyOpttqJGIcsQYfu8
sVTHREDIskYcmRpz3/PHA752+heZF4NelJuicdEEvafDBNGHmG9q2KygDHD/yX3XFQeUHLcmzvG7
axvnHu7Hb5O6nz+QLmOPpBpBcJLme5CqutpCNNttQiKOlMaMhP6LV1sP9+OaCvunuFTXNbxCVv7J
5Qf7P0GaGkOSEwnZiVMuzmOjv6V305OfrgiGF0Zp0coimRiz4kwEJaTvarSQxK2qe5VWAdZGMTd8
zAZTxun1iiFQO6lViZqpJGsdg4bDxKXOVU0BW/ZBh7+F2t2bMciU5hxzCCf+sITXwmv4gF0J5fiC
GOFDP1eTzf8RzeBPgtTE4BsOT4MSbAXRrXwLTzV3DPF9MWnrOVUwPTl9mdLS9ohPIAnnemYK+R+j
cdUrHfORf7ToBM6/WNLod2JKpM4/kEik08/ILrj2L2Ey3Jhye9zHFgJ2YCi4j2jXeXgjmYGRmo3R
mMibCoJBH0A6WFJQ/1hFiDG/YsHt8RfEySW6zkXrhQHl8AW/2LDxIw3qdtOYbfmKgnc9HZ8cnFFU
BChYP86Fz3rYO1kHIw+fPQ/3wu1fSaFi/n6HN1MUjTPgnUt8y/exaw9u8ozEZ+cMIySRbBuvNlcT
FcbE6Q4gLx0oZrBlOkHBg/FUnq4Y90tdZcEf+LW8QhKEu1uVhNjtjZVChvJ5W4znE0gWKULI2gAl
A1trHpemkJesGHo8mabQ/ykrK/+Xe0C1zSZfCEGHJ9OSDOi9sZVsTmEy0uOegH0lmIOnkholV8Ng
YiqrKPPBnwtlZwYYug/faYNOiLyIA/wQCJH/+fTFEopl/GseA3UU9KOT9ZM+DlPd992rL8sa1ZA3
JdN52SheQDph9wA3xaoiBylHPGu1oOpgaf31fazoF4WokSgBjPbNJqVmkNbgzCBpQueeoarM9kYu
ctyg+pXhjkzdiAli+bJcObfolq+oI62RldpFKYH8D69AEbxK229y/ShNeU/VK3JdcyDwyhHSh+Ws
sv3lulky1DBiW3U2SCa0xK1k2FV+OOZVtL+Mq4AxZ9xGL+T3LLOnutBqFh4MTbCGKuiQKIF70qxf
zeKNaeXwLdHMu4mD/KPXHjyU0J2XzjQ73oxoMFEZylk87RYdzPpU3DGX3r2wA4jGmX9TU3aP8tLW
WLz5hXjpg8i9X5wNN2ATr5JtT0IR1tIztsID0nBoZnOe+DBbtmkIkLV520T5aENvOdOhXN3Ttb8R
mNVeOP30wIam1x4xaIXR+js7ygJvkdPFu/Vdr1dd38nbl0RUydOIZqVjYSMMXEfLlEhsPxI8x2g2
7hA0HhcDK1FXABDwQFrx3VAZlF1qg7s0XThv8x/uDkr6HalpxwoARVp1uxmxIEDh5bcglSZlq/jx
VLFhJ9bV+8lEYqZMOMGV+cGY/05BMUT6/08GoNTN3xyXjHWOGCCWisZvddLlqG5iCIiCGcRtiKbV
/S1abJ3ScvCO9gkViqsGtgHZYJo0GN3xM4IXx3Y4rPXKbJUwsN4uQzy9vKM9OwQd1Ir14ZqGiF/N
0gXbt3NiwMFzxi2Re1NsmO6eTDdeOxjkZ3+h5/kkkxDRG0+VW/We38CS4W099slyLgF7WvzoQBL6
swvXPZxQj+Jynf2kzd/Xktf2n+vitHaxRcIqMoLg8QWEVyCts1xziYfLT/7JozbdCf7WCrW6hu0S
FqUNsmq4N6GnMtd0nYhY0i4eW8f8J5bdrC2/kVL8fQcGL3eKjB65sPiQ1DxKogmgZB/admHyBZeY
pyWqQzSKzyEad6Ma6aYSsYaYXvylUvmNxX7SAHX4CmKqxCTKtK4mVRBXJcMAniL5KQp4OWKNA9xt
HTV3sLYWpzv7Dm0s6W+FrUnTkrTsOgtHqNVJKvGX13uiG4vYy7I6Iymu9kHJIMVJLzoqDKeFTrBe
3D/xO68eBqRB4RJnpAS/s/P8MIPC9jA8u7SsProx0KCjSykirI5qimU0muvlBFYhtWURdhSZ+9A4
xj7iDcQ93yBbVld7aB8FPB3FX/clZkssnf+8gPA362WLtnniE3is3nC/UzfTrtC34/2NWDzbWyu0
3DpBk7xxbzMzdhWVCo/jWyjfWZ8syOP9Td9hXEVn9ljQC/2IPIbnMiPW9iU/eYLGxVr6CK/VtP9W
cA2dDY92NhkRNm3CS2grOTW+8hKbaDQ9iJQoxsmGvHKGAHMZSYX+3DsDqHQj2hYU0pb2b4edSFys
rmECAKgy4V9LS3nnSoCdNfrujoYM1zoR2VbJyRA1gv/1TiLEdfkurjDEWpOQA8g6h/1+UIKHM6eZ
3VFThfnU3K9H1FZj8VzehnfmrB3es4Eudw2byuu+3dNPK23R4CotfRtvHi8fuP7xPm5YWGPfO5zL
ucs9qHfXQHO+PtVdURQ3vjJPW1pwg9zREojFNLH8rNR1AP7f74iaFqnTbFe1LOIk4ylQJVTCyCBL
THHnykbe2kw0kz+xfToRW+x0vXT585SbLGViCaUCykR5kxfNWRejV5cfKIXVWOIA3owW7AaE3T+T
czKfCTvnJ1Xr2dD1blspHKkatuajXcxkAMDWpu6+xfJCbYoRJDbS/OX4cNr2CzDkSXF4WNbIMghY
JgCwreDYyd0+FWYG4smh0hRdXsWf0Vr9KVBsoSEV6HbIx6jnY53F0Do8H5QRSsFLUUmUBtdro+x0
4ZmjW4GqnGcBP17ahUJPEGFIqMHpMpuumBtDtbXuZ/EH2Bb2yN0bu8TYk5wqsZEFPqVertFCNjJs
mAgcP2xlLW3LBp0yH7Olepka8uCkJM3BiPuJYm47DSUVDfWfuQW+f6oAgJVP6kBxRFfeI0XpFFSt
JjWjnkF98AF8rqg5SA6ofjUf4xDs0S72BgdwKz3fW+PrhFE2o5NopxZV7PMkw8m3BGzYCDqyuGYG
AB2AscGzGZ562NjZxfW7fHuaW5zTre+VEy4YQbBNAGvJ6iRvgDJtQGcsSgLwUwKMHHPAHvwdl4Qs
bVB1MVjjanKBulMrQ9IX1Pt321Z7KnQuytcHOVXCZg1S1AI6InXVie6GO1qc47dXiV7pSuze51Xj
9oV+Vjf4KF/iLuFkX0ZXg/VekRWjyt84oooy/iMd7Xl5LBAUT07FPyae6k1b1R+ErzY63VuNAQQg
DVe0jIppr1GpY6bGOYlw51R/6WEjwMg6Wa1gq4MDfRr8B/i5BFTq8sVEsd1I//8BsO1hzwgllyrd
AUOLVDA+RD5fbMAivmDwYSRN35UQFH1Tp7xcL/DcESOkQv3oWG4U30BW92W+MwcLipgwgbNhSITB
iKiSwcNH2U6vXmOrhINQW7aw7LSOR2yrAjbJrxkGQvRd4jFs27asMqxCRV1Zi3rEG3ta9YS19NTD
p+S/eNuK80q2ugqsedd4/ZA1HUsLig94Yogip13QeRTLqAE2hmK6bFvC7LY07rnTlj75+h29+BuR
ba4vpSdwxODsr5lhcRJ6vVZrjA4y8Ig4uWJTzqre9UyZY3ILHvzeLnrkWJ8xzBE8H96FxcVRuORR
4kSueQ6gP8w1iamqbQeUMbi+reZPwumz41XAuEwoK44uxXGt56VcYQr+pMTsw7ipYLE9R7Rx0XnP
65527xV8zbc7il84CCokYn7KY3s+upD++9xxOlfkZ4W3hPmSW07rizv0k17BLry5SwJS1c0FvZbT
lg60wSylOSREsaNVjGxeuzVULGArQqypP/oT6wIpMHnEpz1yI+p65XLah61FNmBUwbN9KG7NlanR
tT0UUUqohujMhpOeL6ZlVvVjcZ4S4wCTEJhAVrpJF/SP/tf0CGLq+GsptYiGwnUlHGKG/xR+ODzL
p5muwTGvv1tyWn04neBA6Y4G7zmMgVp2btUK8SIT/n5Zeh6Dsx+5C/dcrc6Vdl7aWFnleUsghyf1
KGfIsBhjuAWZBkt/WbaNOEqrMvMj17vSzH0rfQ4Ipu3OZ4RL5c5JUk199TAWOLMH8q3wOPnerEzV
GPlH0271g18WEpk/Qe1inGR2z1pXeZlheMzK/sYbT3y3H6yWBBw8Dwx2q0QqXl8uBAE7adnG/wkc
d5GR3VYm1Tuu/+gHNXOTf3etDN3nxvA0ychUrIoeq7DdaxbSY7qPHR5fGoAL5p/1nGz1BYlH2aRL
GQgNNj9zihlwIK2t0S6QoBvXuHXMPcIhVqK3NcQkR6mPYweA4vr3FR/lJsOf6gu/fz0kmizoQCt3
DnsEbyuyIlKTHIRpa9j8lyu8YjbyYXQuap6hFpdxvY4ClFK7dlOiJA9fjtfgqa9zvmdAMiJ0g86U
P+JhriXiHEoYY95NN8TzTzXxPa1pd29U3ZO0jECnK2N1sPTyzFFKa97rWT0H6250O9dF/EX18cEn
9MA8C+StyCbEJ5UNYgk3g7HXMnd9uehLXcWdpv5gQAi/y2TK9Z+pXOSkF5+Sm6D9I7i18B9L6M7g
LoQR+scpE5Anv7pY7QoYMwdcf0Co0TSHzv0X/XIoXzuFV0INpgtG7JipOITZ/AFeEulLqGNyvTGi
DCKYICF8zHw1IWIicxBLYA4IsOu7oEkKrHuVXlkeL8+Hf1bjCWSkClOxUeonMTSUNKTsR1FFYnP7
14/l2BHxlrVogF//+KKdZf5zFvJE/m6GkIAAZRE6iHrYJ/J507cHqYmLMHskhA3tlktmaIo9VlzQ
88cvaPIJSuQkne5mVDLGbiSuXhhScWLvo2v4/uzxS3i/1qqnhRU2NAU1JCG9On64A+LZcOOaK3G6
Jo8SAUQ6zVdD9cxKbZ338KyH/JtIO83G15sIt+2CBLIgLk27isBMiTHmURoAa9OE8068Q3Jaqk8f
kAJzeMPUDu84NaTSAnaPhxR/tjLC9EElTr0O5l6by3yzME2kWkaAM2Q3/2Jk/8D81BGw6ifi5oZf
d+cp2Doa6yprJb1GC2w0tQZL0m6krTvPYISO50KjGXPWJ389YDJAn5Hi6hUT8jta2NHHwtNYr0i/
5hGnLlOe3sYF4JKcE17me9SpgbHmwYJ6+srnI2/g4Fk5gUtMit7VhEj/tixUav12F1Dx6GVGWNqn
mMXN/jtjMkv6UXttln6+MyE15Dojnc6ILQx6f4lkM7PSz2/eKgnAAisXToQHdWC9m9jlKP177674
qhuSM+2JiudGU6TjMsDHl4c4AJcg5WCkgmNaiSwu2KxkES2Keenwm2xC3Hdiemp6OFsFs+oMiYSC
XvLpNPxlQvBzEXKAl1p7XhQAWIpnF4L6RqTXTrTZWKvJxKzAI9EPThidzr2UU3BM6l2rcWmunYLN
oj3Bh6R3tuvQBt8WjAz+NJ3p/oqiBbgj+5r6uftwK7MrSg308dpX1DY4AEJmEaIOvVkQCgbS7KtL
Zn1pHA+uNwW0qojKKPkQK41upalLCjCm8omogka+da/GZHoluLrjf91zGdEjz7PgSKjp05PlgbAU
qv/G0jcL+AiEtE+TXE9yFis9JjhcG7sRrQPIyRP/HBj6ufnzyoI5cmjtWRnU/oqMouCxqIp4gayf
2OSUHIHyGgEVAyHpdomN4HpTBo3612XomzcqyLdhZlpo6bte4qANbaPdstUMGKZwlQSt2rWCpKJz
eHNgGEDCIWZ2mybg0Zt6uTKBSwA0LsL0c7qm68qXCS4baW0FxK8LgoV9nHBJKTZtcl1/hHd306m+
3O4ZxlMff5Kge2mh2N4RkeQOi1TAXPHb4t3EHTFmczk73hCRwoGYM0RhJVSYUYsszL083ZUopPVF
EnGzS4K0Zj6VCro5YURK3PJ7yamzzd02NqWe/Cm9gvpJrHJ/Fj+LVZpsqqkhOuuEOLMip7xl3iH0
sG8eS7/KUqTrTnZFiFxSXNaMlpWDi23KHmb9rfPCc5yj2CX9hEyvBe6VimTqQc8Hq8SIRzaPajlN
4cmIQGgXjXdSxhANrBzq9Oht/uy+iKMuFfmDptpXlaV9znYxEyyNLVLnqxfcysg7Hxl9F5+BdqY4
zOaZEWH9K6atH2I1UT9rA2xpmuAKPjMKxP4l4Ua4+UJZYoW5EsUK01jZB0ukEMFdOObvOo0LlKlU
9iqa5RJEgtgUKfeQeidbBjwKeY0iAXTwvtCS4m0ffS7aCGplkOJvmMA92bUzxnd2Yh4HUmW9HGE7
OnjCXi4p+RZszUEkVn8Hj9aUymoNVn+c4UbMnyr+Eg+/6yIlFbIg7JG0QHvjz2/d0GOw/D/zHARX
AnsV87oHE1q/kcjMxv/da+vKMIFcQo5mfDSQknaE9OJrYa20zx8j+akkco25GyuKN4vpXGu5/WEc
0BM/qeLAz5k2BULJKySu+SaY5XnjWAR3gbmRoNvRqqA1nv4lcWxXR/SDXQoOBPXqPb/72MbnHCms
AAYbInx0gaY6nqVcf/vJzmL8BwOHOVaxrzsyHTKP15nw8rYHY6Du+zrxY8QhZDKA0/VCVR2X3uHd
Y//Sw7rkpic06mgVuAC7H0j6THbeYE3evCkXTG9yiLWwdKaeMOv12+08R+DWnBAB+SK3XLAxW2h9
1wjv0No0/lE3qrV19cbw6/1xGf5ijh8xS8/h70JRtlv6EVBUDDb27Rnesm0c1UKvl8fjqRDQleDz
w+IRLdlCDZFcgbHG5IfOrPr+ft0LZyiGguHzMxn7EjS3lE6nzIVJUIcRdP6zfrdMkAdnb18+awEr
WCY7D7aUfxXgQ1aRUwvpxxP7yJmkI/Gil7HhTm3OnSDtdgJeqPEUmRyZzFjDAKEeUKXs9Qb8LF8I
Bs2CCHW5EPdCP5OoEhQ5xtDp1Vs064XGbNh+z/3yKgDN71ij9RW0kl1ZjTgRa6qYMYim7Et5rRiA
pi9jpRr/f7h7kcG7s+wbGVnVj7WNf6tlHadDJr9+3t+MThvtkFkc29+kBl4//dQ9RXxPW9ZXCUbN
qC0T1Wnb0lS0KItP0cMp+JCR22odx7GMRsHU2c+C1GTsbIgbhvBUBvyws0cqula4CrNcE6IYEcKT
onSCoIsOiMqgjgH0KonK8evtgyViZT8uN6sFkJ9ItyjE7cSLBfFiLTsJBtS42x7y0gkEvuB9uCsh
xkfpggCAGrwgnqxj1aPHT0/Ao1pZkFIJIQ8KTh60FLk6tKtlK9k8GqjPRTNM3GWzJWQd0ElH6Di/
tLcdviznfZ4jXk+nh1T5iZpRVT88MMMD57DosEIeP3i1JAb2AVtu1kJVQhmcTEZiPFAuoCn5OifA
iJp5uMMBgOp0LxtME7hZN95qJmJ7wjVrkq/W9IKgekW0jbj3+FUmgIw1ZxsnhzoFvLg5sZ+V0FmZ
ncbzRIziFpDaXNvCHpaSHEcjyruyZUi0H6GwqcFvUBUM/X+ctBNAs+iu5RF4k15cFIAEuLpitJe2
O08IOmwjpa495yFHsUdsSLb4L5E+p7HaHioGphD+jJs24JFho5obcPzAlbPOeJFJx53qbpTG3e+o
GocHFcNSTrNWEmfn3MAUMQ83S0OkygiX/Ac7dfHAB18MxkLwA7MJ2IBbbPJFTZSx4OvuZXrLXdn7
NRyN9qhzMQZWEFUFz6xhZA10Z5piJyxF2vIU+ba8QznlZGVIjkLwWv8HfzznFrF4aJT90IjD5NXI
HOLlk5AS1IYVFYaAgdvbMEs9hKkEFefwYo8+iOUGRhHwBxXNd7MySKgrgyf7KptjThpNWFq2ybxY
3gdObSscUD+ePdhBCnUSstiWHLIeLfXRgoU4RQ8ilOyGOzOdaRbYHLyCvCt/3nB80CL/XcUbEuPE
Q5QGu25PJSq1Zd2F3bur+FEFXNug7N7+R984JJ+U2PNBwVsAhYo9Zv+GGRnwcx16sHrEtq9sl8Jq
Kdxz+CEEAVDeSkhOi2qjK2/30L6cd0mf8pE1MNJhLCuIuZGtLwWK/srwfdBDF5hZSdaScLu7ss5K
Dfv9j9EOcw4gzN6QgwB7IYrlQxMUUVePEYKEk76j42242D/kepQs6t33XRH/UGpEtyYCnXB/+ZS5
S3zMZ4HWrUzsDe6Y7HCI5twAUQCx1ceBlNyUCr9Hu4sQStEK2DKy4K1IXscQc+J/d9WkJVG+HXUZ
xb+UM8cwgF12W14Tjikjt8HGLQKDkh0eGcS3bm6rROE6Qz2BUPxcSiVBYKsNMyDEYQyAsorDIp0s
9NXseaCUZGasyd+zA6SQe9EeSbqO9O65N0zEhEu7umfTuZ52IVrtalzxVe2ULpvPqfDHx+d918jl
ebQBMq0EqQxWhJa3S99iWC+HzHQWiUaISUNXLCkeZdJm7h/8eYNHGCdzSmVzgytoh4UUaea/Gz9r
kQJJxhmhmC/nQ1wE/UK/qkKMLbrEXLP7nvhK8g73f+ouQl9sMkwA3lkK8BA5YG1lqUUcUfPquMai
1nMhwJEjD94k3HB/JH34bWQJ0EOgOAYYJll9jYLkMJGRN3ZiymeHB1M2WsNUPn+Wq4uwfYE0BdPg
+hR1xpPwfGDEMiGkNTXLLAFGQG9oPae/+ruaxVZ+nklaDq29I+RLfKxtZOvzMJstiGNHniAfS5Kx
jSEySATjtShi9fA/6BZiFnrSE15Y3bguXe0SywuLg2/ufGw9VPfqnvjZKRClmVecVvdxYu69Ztxk
3jvHmMCKkyB2UZLeBB/WhV9Jz88YpsQ/UQSuLNrnYqx4otrucJfbUjUKictPNilWZp1MjPd546v9
lyFOOhsYvCCln+GCtvXgDuBzz8UN4d0tHw1HMDLWwgYlYlMyF9tSYA5tSGiGNWpUeqsy4Iidj+19
+0j6VIgaLcK1vAdQw+jvw5L2lQ93OKk3yfirAbGNwz2esjuXwlO0vH+Z6QD6sDTOO9KZwCdVzGG+
7wfQ6RfHCfU+aYDybWNTF90GzCo2pAMM8A0R/x+Bki9b1L9+9sRhCGQ8BgRjNvnnA0Yn86Yz/dzB
SuCifKe5EcaZlG3DdGRnVzbjRA5Y7Jl3hx//xG4+MhAeUP3W5kWN2y49/BHdv8HqZeM12PBp7YOD
DqAHFsRSth+Ifznx3vcoIoH0EHlXwoV/V/hvzxtpFmTwG1cnEF+Yz7MHTkem/gByGuqrYsx87JJZ
ukLQbMNCEyw507UdBlbOM4iBQ9J+TxGKMbwV/IjF7kGYlMxeUH4Vb3cKEZcCltg6vJwjoybFTIt5
J/B/CJCJV2AoACJCNDksn9KoOWeHZUnKeIylmKcKTaaU5sP2sbFIZf8mxYkRHNhXpdzikZU8hbA+
yErSa/Qp2NlfvyAh7oxGnYc+1ymaci0zmcuAI94fn+7kY4NoHaSbuLUb5SqUJs5U8Gk7vf9CiHdw
/ebC3VpA1pmJvPIZuiFsK55n+9cclXijT/OxclmmErY2Xzl5PQ0u9ep3m9AEjwj+sDyoDO2wXEFt
TOHjEWg4fRq56ITTijmZwDGdxp4ajGVkROkdzkphheWj1YjHFUwpqK+InvLdAcaYl9LWyF8X36/g
yMHDHJawfMnA6xUqJni2zrg/oWYszeOA6gpvZXD1VfG77p2YPebdTKdh2UXGBjK9poTXzhf4tBIk
rVtMucv9gTuipVXGuVTsAF76ETWjzombGOJHYcMEqVPL1Qb8P0WatWY0Jk1tmYsaJVXVp96SZ/kh
VvIQVuN7OVt4f5GLX+v3VIhxgdwbtiWpZV5cHiFmYJTWWEN/gSaiNjKXLY1jKLnubYGYr8r3X38C
tHGQo2nPoV4ij+MfLg5UkZ25qcmUKksi/QPMpR8phjhzm+XagLTLusVnQ8b5+qNG7MF933IzanEb
e0K20hq+i5dUvyzlSckYPbqhJ2YQM8l25M2BtXPMHeZLVzYwrHxAE0k/AGdei7tvldQdA4UcEobQ
bw+viymbMUhxroD52UwhG9cUC2xE+aSNE6P+wTeHo2NMDHGapatRlZjiECJnHZB2zANf8T29sHvo
0w+hHPjhMMqVJEgkV1WYE2U8qxhvgWFkCscdU9QicDJQ38J2wJKZlIIUWIgqwgZaxiyYaCCoKmzo
aPBIGexyJQz7vWVm1v5rokXW6dzYqizWktyfHxujydCF05ChSKKcUQV44Jm3pvH3b9omNEPARlSv
SE661yHnKKdBx3t76aMo3xzTq+tMEPchaRK/EiaIhx5Is/2RGniLKRhuJQYMGjx+f9QVKiLcECUd
84er/f01lcaYjZGocJbrlF0/YwkbvUNe4kB1x119lZhLVs26PCI/LvyTUjSV2EtiJiKJdRvGUXUE
vOHijpL43h/kKzdnXeZyFRHX0x0pM7PMTlbu2iV14yyca2PLaEQuFR6uZv3soF2Rk6EGVOB1ajX9
0tE+ry99Vd7As6E2jZ0E+aJxtbBfrTnpjQMKg/5NItxrU/OU3z529+ErR7FDjFNEi5DqcZQyfIm1
yGa+Lo1k2TIsIorSb/dj24Rj99v8VsV9+OWE4uDHhGvsz7XYjHBrWOhx1qcrCApn0tF3IgFZZf1n
IaTX18MjkdDLIB20f2+d6/0xgGgHCWGqZEFORBf7SLFEWGBzVig0Uj58fGxe2+td2vbyrVDqY4rY
u9KckSyuWuKh2CnmG/CfUeV7M2/5ybkn5hltaSx+hqzxzuWCoxa3/88CRQGZK7eFOWneUMc1YGNU
MAlitYHtmpxX2AnB5JCL2wfgmLIVLe3sdwJ3RqxL7PNH5jk7kuIUljhWUCf7eS1rjuLQ4cAdLAhx
kqGqqG4OEKlhOAJn485TM6LARfHkrRglwL72QVPzNM+SKqJItvnsUBZUgw6+CAexuL5lXgryTblh
T9RD/dVyjXIO/AnV/Bpe74ixk3iG8IsHqrVU87lA7hU7kaGivbExKZ2vA6nuc9AO/7356qKMtose
mV83hN6vjmScYDFG6PJcwL5YbX2ZfxXYZTwQd1rZxubBIQMM1a3Q0EDTlHxaS/VDGwHhz4GIzB8j
CDY9vWqd2h/OBW3uIyrgiwlXYcf57owlQ3+qQQ27CLNcaDDym6S6WJ3+86c4HpBLpxK+cG34Aahk
xfxvheXUgkEzbasue3GgYKcnHFTk8uZa6GyojE5rx7U/Vd9YUylhEZI6Rbx9bcsEwqM2Qq/USWwZ
ImGnIlsNX5I8rLG9pkVFScEJZyOaUwyyIvLyEE37VbJKPAMbUzwGo3OiF0faRPkGTfuctTJQMPH4
9bQGfGwsOM/ArKAZ7/vAXn1c8H0Zicuzxsx5j2H0t6/iLjcFjTjceh56W5jD2mzwqWqETKHI/zrb
KLKYQu/dy5Z9O5rEJSBW78cb9SEsydpyDInxsAdDVFyeOYc4ri7kgQlgXjxFoEAd4CPJU87zw8pR
r/7+xQCv7oqyfAI21pZuuZcoK/AYQF5kwgReTqJQgdSkYE1fE/7FaZH50NIvsvLtUDWcr39uSeeg
qrHxbEKM3K4D1mozzysFelD6+kBExP/DOv9ReJLEFkL7ligDsW8INCdAk135a+OumB83x6DaljYi
ow3AXKPWbdRblod6oDasBta/M/no+ofi+9uk7a5PUj2Hwxv7EP0LZ8vwOrIGKr7Fa/hT8Ost5iLi
9FDUzPOUiRD4HarhMA0HCriATQwBDiYNK6ttEg9Van5RUaq7V9opcSCfGni33wx7jlWqtPrxfj/K
YblpdM29yIvbTBk1aQkv67fyJMRT+H6UAO1unzNQ2x3Rb/6xll2IO/KLfW7+WqY96wGODValqogA
aRi9vW2M56JSIXVUVjCnxiU4tGsNrg7TqJY9vCdz+KGiy2Qd+7t31KmVlIe0HFBk5q/hbgNuk8w0
yla5s6BhJJ7Y11lC8qiY6Bdtk3GTB4h3JCLvatNLHDrpIRaexx9iMPlFr5oZXpYCVEUOUiifjrRt
AuiHxkQB3QTDKN+76xi3OI6poK/4o+pfxiIKJakbLG6rFpEUke19ZMDtuE/uQs8o/0optTokGA3q
/6DB8G5lS0hxiLeHnbc6H/lARO9CExCKx9c1rxYQpHLDZfs5+RmpEm4jjVT5t3er7+6TjO++SXlN
boCdwFywOdWOCtilztj2BYOkaMxh6M251uI0dAeWenRIxRlneM8w3+TRoyxPGDUjsEgbcQjoLja6
oTr39mS9DWpRfaAu45yGR6zXeWXIVnH0rWm7uQ9TrWeuJEUKtcBRAcIY1kNGbH0WN/1pXQbXDl3G
OmL5eCvDNaePlPm5b5ckXD5KjFZRedIntSniwh33ZyCS1EhM1DwgqTTxkrpBazP0JYf9C8/bpAdn
V67l4VHSL8oA4pjSMlB/clCReZLpW8qKCsY2JUSJKwUxh1SO4RTB88UbkrsH2LDdr+14c2x2eXs+
5Ii5fFEeegcltydk48wJE+VKRrZKYDi8lh8oAL3D4NFgFg+va7qJj+naLRMi9ET8Barrlef3H6kU
3BTAjsOFNGNCfJMQLgs666ACXYWX6R2WL7an3EBhP75r6LZoXYHzUZJ6FyEpUStV7RJxIvoYAOMW
ESOwd9BXXQEb+sijw0JSoIXooKUjkH+zC/5O0QYFVR5LlfFWVOyzfIdNdfq/gLq7YU1+pTX/lBCp
fuDESCzhBnm2UpGvyfS65hixE+DO0Sac5mwMFePhIzMrLAh6tl/14/qTb99KE8+m0F7jI8czHZLi
P5JETWp/0lhD7hiliTOTjEcSzXeBXpGZGEVtr7YfYnGuFF4pBtTPdc6Ls1LFd0+kyprbEgPZ72QZ
F0kh8a5C8pOBZQiqXoNtmrrmbhc4oFGPSrRh3BuVrKync6GF3P2ANKkZN/IPE44aGHe/wGWWhVKn
fsZIKek7zUekB8coPzImD5DWlioZGwMzKIFDFBATOpruXWi4nz67TINe5XQFtKLNpug/55OBFk3r
0/ckdY7LfLLmChZavNCKDae5yKo2hq7XcnFApIQpljiqN1QkOj4cR5xszxeZTwx+84KALODNiy52
kZoPZoz+hNiMHodEhYa2qv3z8E/cXdbUHp3XXCNShYJRXxx533oK9WquGu7vcAetcCAKsMnGZiaE
GmAuJLMgoxjrTno/v8FW3kLJPzBE2AIBPzDP46TRVaWmVqok453xzEhHWZjNVWW4lLDNQlGXBRSd
UOTZfCAzw794lAWwNCFgC2Gw/DgJkQjGVA+AZd/71kZLMrzP1hToxbYaS7NFUTcdbsyMbfrFVmLA
SNibA0rTRu8vNnoBdKB8XRfguUgdnDrRHCmmo/KPeMFYvaqQuFcMGXOu1Wrf6DYjCw/UcC4N0fya
OKDe8R+g4GuDrNgsXwuxK/VLfpUPmoZL/dXFiA4z5isgXXJ3E4HIje9mHd+YR/R0RCmgHjrbgY14
alhXGVrR7tMyPnHBbIVyvYYbn6jlsHkdrW/ltsLYs79hHFEdQ3T4dj78gVNTkJ16n6iiztoJ/QHo
EhAe0j5ZLlfdVvFwVCNpwN6Xe683HR9L+D2LQoY+PFijA/5O8UcAkdsavhwed/qvQXUV1nRgv8Sz
LGjGDgFcAiJRaVT8e0A/gd4h34LW
`protect end_protected
