��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����,�1	�)��&��(��H����dP7ɨ���:��0����,�6m���Ib� ��JK�yUh^��9���E`���K�
��Q/��V��T�"���-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_d
�t!���N�S��گ/�TNM{�C�5���M��;����L�S�:�{���\p<��)�0W��B�R<Qt��Ԁj,3Ӂ�v��`s�HW��眣�U�Z.͓k���ŏ�^�sGt��P3U����ŷ��T�ŋ'�Mz�w��� R����]=�0��=�1��Qz�Tl6�Q�5 [[̠�H��P)�x �>D�XTV�fP�Wx��bNCO8X"+��v�Dz�l��Z����h��]�ūoÙ (~P� ﲵ_r�N��@=r/�D-[SNG��u��(���R�.l��`���E�:;�]���.]ш�(�(z�KT@{+�;��0Ne�����B�<�z)�����,���ݑ�!a���B'@#�l�Vϧ�^�z�0���U�RU�a�d��a@uu�M���r�_�%C���b��d|���~��!x�9	��¢(�W��j@��E(�>e��w'���B�޷`G��� ��% �åB>'̖��"� ��%%;C�e���-�l��Y
w�%V
�H�f���8�\4���t��<�m=��\Ey���M*� ,ȩ(���T�[���m��5!���{��2����tz�����K;ZB���Bk.z�>O��(IE/G�h�u��j�����`+*�����t5�5�+�"�dA��K��B���,�M2�w��,���B�|"���s�"������)"��?FydQy,���%H~����7P� #�]��tr~�n!�`�bH*1�P��%��wl(�R�ؓI��T��H�?���4*�I��١b>a��{���g���N�WxDR8��OZPGź�
$o9�c{~�zSʜ%G��T��o�˻�� Uj�m<��Y�m��^�w#v���|�9�h;� 7�ó'R��O���W��|�=A��׹�v�	�ǟ���e��5�]Ja��K3V�l���[k��K�\oRT����C�v�} u�!tP�)ȏW����J�(JX�lbU��15�*�[�[�	,�>�#�x�9�j+���HEc	���w���0{��d�Tg��Nl(����_��}��p8��@�42��).��q4ۯ��U�����9��iyZ4��2};�S���v㾓���$1�oЎ�זũ�d6��W��Sg^w��NUȥ2]̄�;/��0&��E�g��Uر�� C���S�l�����g���s���&g�X���&y�o��pF���c8�T�g�
��
YMuS�<�[�OL�bZA�4N1�J\��\� k&T����|A�`���8Ơ�Kn��SնS�nk��6���M�|�����e�v���D�;������'R׸��p�}PTMP��ں�|=���o�⁺A�L��,�N�$q�tQ���c*vh��������j((�2~�a�@C���׬h���ʣ�bD���4F�H��1q�#�jC#N��e�0���~��2����c��/!/�[�[�U�O���G�������D��l�[�+{�'][�	I��4Dԙu�q!8�5��Ojv�g)�ng�<G��wCX~%�(�-�fFK�޷v�Թ�}��K(Oɧ����\��.⬾GM^�k��ܓ�-G?'��w��0� ��Ζn%:��' Hї]S]�lΐ�&ν�ܐ͈N��<���8�6��D�J����L�a����$��S�>��R��h�w�#��V���"�wx�e���zr�|t��{
�&��>Ձ�*	PX�ӓi-�I��R�N�~��LA�V�{��y��������y��M�ܛ����r����08���;�O�b�sW��!�@<7�dk�3/\8rϾ���_<��d���V.�In�&�L>��־`���'�S�Ti�k��CV��&��S�z����~�yb�KS6�@��M�8㬓H>�,��<y�.1�W�P^*�K���&PpR�ay0��ə����;�F>ӽ�(�������P�zX0��rc,δ���\$�d���U�����3H��0ƪ�)�W2D{@+�&t�D�����Y��U�.���:a�m֠�k#�áL�겧�."��>,(%�E9M��_!D2����sj-� �y�����a߆u���!�_n؎���9����bי��o����,�W+�]m�}��n6����6�{+Ҙ��ќ>=� �R�QB�+���_ܬ%y�P���$�)��g.Z�L�~�|��r�����2|B�ʭ�M�''��A!��C�g%&���4_�f6ĭ&��^\9BQk6.�P�����;��v����-�8��B>1J� ���yc�j4.�6/��=�Bn]�A�|�+���4�`��fϠJ73�) {+%�;a�#uM�es�bo.D�l�<�IT��{�I�ZU`����iU�Mq���5V����D4�7;Zp����^1̱��w3@{}۸�Cf�DyFcA�I�79a0�7�^j�L����3ӄOʩm+���3�5'2j����z�;0�Ї`���2���R������'m�Gߨu
�`X��xj��1B�7��]8�Oڰ�hkB����Z�v����xg���h��"$��U\) -U��b��]��ùy���{"���^6�|&4�}�"�2�$?�Nwd�k /���j���WԆ4w�C� c��V��S\����@O+޸bCʆ�:���M��~�"\���3?���mZ���-�4�4�d�8'!�i"J���o��{*Unl���E���G���zZ����~�MԂ�5mTұΠb�ɤ�	��e)¸�X�_�Me�F��Դ%�b2�et�����<|�эf(;�`�I�k�>���a�eB$� ����|B5Gn�zg����j]��Q�rĩ,�ϚUů��ҚƮuwML�2�W���aQ�KZgj�D�p!h����Z�m��o���]Uضd�$m�C�|��J΁��D���j��7d)1:0�V,��袠
:�Oф�m7
O<�6P��}�=�"��N�,}A��7�L
� ���i+�M�P����|�+���;�<���u�7�����a]V��bU�P�1�|�9�uą���}\"�?��j'������L�P%?���w����ּ�ϽO����q�}�����~���ȥyc��ߓ���vZ�|�72�=�� �tC�䚯J�K��E�X:�����k�R�
��� �\Xi�b���e$Jy�6�n�sNR�+:�hB|��I (~QI��jQ�m�޹��5�eʹJȴP�3pK���m]������(���&y���J���b��D���3�jI��'�zW�Fܖ��;.��5��d�	gAh�����@�b�5Rzb��_�C� �!�`���r���x��T���ʎ�7:T2���H��[v�5)�lq�]}�
]!�ۉ �ʸ�逢�%R�v�������Z���լ��;�@7����/��b('�~@)@�%��th��p[N�BM�G�#UE���)|�8�����+�f�zՑ���p�5].���E�26>�w=La*���H��Ȯ!�繲�n�T�����R.>(/�"��+O$U�-XS�l_��-<߉���c�M"F����?G4���B��?�2���G��ş6BL|���M��z�����[�r(d/��M��~�证�,D������~?�ң�c����\�{�n�I �y�^H5�2�PRs�ׂ���eP����򤎩��h��ҀL�G��֌��22	���V ��T�WYYb��+�b�ޗ"�Pk��
��.�"����d��D���|��/LZq"���0�?ľ���EX�3m^�^,�I������	P�I�%*?�d�"�S��i��l�ӳ�o^ǥ�2k���Ԭr�a���A��1�$�0�/�k�Lݲ'CBY�t��Y���\�a(4��E�_���tF\�񘟇%��w�GA���lix<}H�C������ե�g��F�n(5sWY���N�pEHU�*>��p	�i�o�/`wK�H7/fo�!�[/p
���@��b�@�0���v�n�W�+�N�w���qԜ�9"`f�m,U_�%�eu5�W�2Vk�n`2��q=��w�&���M���ё}��x��wP��C�7|9�
Α�c�'����e6\L`�Ξ3}x�e�Xc�:�K���eb�Iv���K�(G!�?����`%W��H� ��R�\6~��z��@t����rG��1�7\$��O��w�j�����ZN��p)����pb:����e�bzᅞR�Mq�����/>@�4B1�����1"!<�sp�n�Î�8��{�c��s|@p�D�&���g. ��̫{v�TJ|b�QA�#����)K��q��5�AlK��j�)�>=���"`��|��B��(���E�?^��o�y"vR��i� �����,x�xXT�`9��?�����
+�A��9)�)R�:Z��ޱy�#h	��='NtRa�j�3�r��aю��Fo���"�~;��]0�m;u���u�l�q;DB�%]P
A��G3*/�޲����{��fӍ��<��U�z9/�� �r�8ɽ��Uڤ.�[��w鳿ϒ	.�Iҗ�J�/Ymtp���_�!�:��Xo���Lw�B�F�����J�%�������Yk-�9�w�D���1�x崴��i�V�!�qA��5B�H{W��K:�+�*Eto��	�ѳ�ě���Ĵ�;?~S��9`L��4��&GA	ՙ9'C����c����j�nޗ@�l�}�C�=*�hDQ�c��u���N�Y�RӏO���q��8k���a'eNp����y�{ެI�LE��UL�ϕ1�F�i�\���I��˕<�3[ߋ�S���l!?~E���i<����gY����ܧ讥M������V�q���9B�+��b�%��$_��;4��j%�`�kg �}�s):��(;T�V}�;�Ok�%��%�C��������OT�ֆ&�л�MIem?MaZp����[(�]�ܳ�u�|����<��O��K�#�/a��Z���I�+�����i5��%9� $,#��NY��][5,����R�_��Eb��f�ؽ�:w��?WpVg�Ǆ���{��$bi�{�Nj����?�b� �m��i_D�>��n5�x[��R
&���N�y1���߂/��G���B��. eb�Պ�MX �I�j17'�'z�WR�	��"J��+��\3��2^u#@�on�|��)�n��)��v#}~8xK�C/7�+/�w����Y]�"�U��]2;�~�+�J3�$����F�?Z}2	-�`��x�x���%z�����R�蟷\�Q����Fv﯈�A��lu�Aֺ~�b��~���C;��}���vh<"YiY;�'c�[�W'�<�y8�㪵�;p�y.�[�����k�v�;��hƴp�Wjl?��|i�
���yы䩑6j�(0�[���8�v��U�cO
�Q�5��㳾��~ ������~=���؍l���~��P:N�S��uW��	o���#��\� ��vs��y%�+�O9,%6H�j9N>��P���^��aT���NDn��BE5Ě�4|�&6�|�{,�y6:e�s����GlY��L���/Y��L2m9�jT�u[Rj�X��K��w��P^�g�hcE/ȃ�q���Ih��J�$7�����@/!q�}����R�u}!C�*���dF(*�~Tܤ����K��(�r�6�A�X6��N��I��GA�V���d%�W8�ucDG䉐;�r��zLGR�U�	�v��j�;�Ll�qFū���&_�3�ǌ���ھ7�	&z{U�`��L}1���B�dU���ݟ��R`�d�+��=�ݢ����;��S�8�7��&���E%1�������)t�H]R�kT���#%@>\K~b�0�\>z�K'D�=�A.v��*�S38p�j���������q�m@O�%�_�:s�Y�����&��%�"���h�V������Sn�����Mj}��N9�\/�` Uyu���l�$r��d��ۗtZ����V��4#}<���d=��~�<)���;w�����c-� %����j%����V�K�fn��c�,P�TRu���HG�a�1�U{��Q��/�\�$���	AM��~ó�㍗,�v��إ�d;��F����
Bn/��j�gS_;�'�䲿h�ֻ����j�iPQz�>�z��l��'V�3���w,�L�ho�>Q�8�JIN<��I�!�sO�i��@���BX�ώo��n ��Z�!���FjZXZ>���1f� s��uv���5��$f����?ް��Go�2�7��AO���<��U�v����ru�
��Q�m���$ #�4ftBJtݡ�*��"�,�-�QE6�ʑt[F��4�n�.�0�1�Y��w�qEk�o_V���v,���<^�$���&~��nI_� I��z��6�*U4%��+KSvk��]�U���^>[<NaKĿc�|�z�n]L��ݦaHG��k��8^_��P�
qK��({Fe��CS�,�]
�'��
�Q���/W�T�6���Ʈ��Gw���$��,f0_~��pt�ۦß?�"{��
郧�=��:�m�u��T쟮���gzO%[���(q�It�O�����MFl�i$���!�BĨ��:tR�'�j�
��%��h��z���ey��%G�-��CȰ[�O��1�<�k�1Ǳ����pS�E�o�8lqƦ�	�*ӽ9�z��Lգڦ�{��T�!ɕ
��yf��/�d���V�Y�YN��.S* _b��_j?��!��F)�ٖ�r|��̳ۖ)����9j��S�8!�S��R؂��OR��tq���+��н��i'z���|���?�*wN�9���g]bNx�D��P�l�m�5I��Pa�f�/0^	r;����Yԫ�eU@Gg8����|���mc�Mn'��� M�������[e�:���Ψƙ�{Y�Sɍ��,�u�
H�&8�zmM��!�Dv@E�hInBU�Wo�j�d�13ǭ��N3g��p�ش����L�.�Õ=ÓHn�[��q�q��Kif���\����B;�p
�W�_�{~������V�0X�y�L�4Kz�)9���0�D8k ]7Q筙*D`�s�̊�ׂ�Y��w��<�*{���eA��w�M��O٠���C�/E�'V[���b�`նɽF=�b��A[A��]����"!���P1��/}���ш�0�Ώ|����^��qE�&��N)i�!,؛@M�b��x�T�`{|O�t&��õJ	�L�PM��`\����@�i���rt�@��xS�8sy�g?�WE�S���/F��Q�|�ql����%>����o�T���D�_"L���;�*n�ۻ=vu�k���Ʀ�
:�e����d�a:��h�"d(+�4r�c`��+�E�!���M��Ր�I#�w�p�f	�c!�h�(�uz �Ò�F�Ẍ́�7Gx������Ƽ�r�y�/��c]��1e�N�5�M��V��[���Hq�zʒ�̳s鍞�=͸ݰ�	���B�_��$���X���q���qqN;c��G�|X#4�4�:l�f��N�UF�Z�ܲ����l�b#.и�t�������%%�d�����\���}H�W}k�c�9ɻ������F@��]
}׿�a��⁾ ��I��ד]?B���� ����2P�=](`֝�jui8Q7R�$}��^Cc�t���:W{�:U�����g��k�4za��g��u{v���AL�&�̌i%T��g������6wJ�'�Ksg��T�8N2����-k&U���\�C~N�!���I�Ք�1w��P���O(��0B���慠��[2�������<4B��)~;մ�x*p�sMrz�m�rlU��/9EAG3�θv6F��65F+���F�G�8���E~D��]���.�Vd�i��(ɷ(>��<��Hh�O�L}�܁4$�9\h�䗑">]��~Ka#
<c�!d�Y�h�9��zd|ɰ���i��ji�����}W�m��{� b�@�����n$?�'��C�PC%Q��mj��a��t?��#j��|���:*e�ı���3�� �79���A�Ɖ[Pf>��x&���,�AUO`����&�+.R�<$�p@�1.��d���Q���(���J_N�x�ٓ�4�����A�2���zN 9�`Y(�3�]"�).�̐țx�p���r������ɖ�S�+rD�(�t���01��Rb C��a��>��X��V͌Q6��`�ZI���P}r��PfFۨwa`�qL�h��G��|���[�n��]6V�15"�b�i�-� ��.\��T��Q�ӓ7����l |�v�\
c(�2�\!���w{�%H{ib��>R�V>��5cE2Yo����o��iZ'xΐeP;+oZB'��m�Wv��}t!R?sѢ�e�]l�0�J�\2,�W��^��[���#�Ȿ�,E�%�I��)����Nm����S�W�� /{���-�Ϫ��\�U�B�DF��O,W,ߥu�z���s�	s�Uq����<'�LKyM�C���8�����'���uR,�a��Z�����R/ޞ��l9������ݖij��qF,g����%k�z�i�Y�:w��M$�n6#��Q,ߡN���_��N�Fj	�?�ʋ�U�"�C��(<�ȣ��#�<H��\��P�Y����$���=��W�-���'��96�+]���ς�G��@��^f(�恾�̣L��`pot�k�ܱuots�\'���#��!�L1�Ц%���j:n<�>�(洸e����|�����(��v*R��s�Ok��iVcRUۻm��l��ʋ�!>|l��>�D_����0���S:��8�Z&Ò1W�0;C=�,z�pŵ��,��$
n;+Tz�mK"�y��W�T^�\~��G(Kk�6d��`�T��:��L�[Yʹp9����yd�E�:mY���4wk�����O��@��a,Ů�o�������<�߮3���+�	�S�8,��z{���y+��=]J�;�o����m\��e��Ԥ�ˇȩ�r�4 �De�.V0�ת������+� ����s~%m��G��i˓�d���N�/��ڍ��@(�ޢ�솘�iIGEb��01#&���V�r�����m�O(��}��8X�.�Q�6�;�AT�=+�,�53
���x�� Q��壩�dA��������V�U���4s�{�c�=jJ����+�f��ч��c	��L��t7�[-|�8V���}�a��8���z�K�`46v�ܧ4"�ڭ�:�����<�+����1�cmul�l���O.�r��]<ᙊ�0ֻ�����=	QS���	b��K�i�����}	�$ɿ�f��M#�ϛ)�S-���W��o�y�0.��eukY��iq���P��,���'�+�b�M̼�v�ˑ�H�4]/9�<�o_��آ f�Y|aZ�$~�U�`Q_�l
5]ݸ�.!�k��d_�*�xQm:i9�v��+���i�-Y�<s_8���k�kQ��f�#��{2��y,S���#���]w��H��/�z(L|�"-@����ڌ�U2���}>r�'���P��`F��^���X8�T��fY_9�)��ĴN��$d9H�|�t�uKA5&��?���������#��o%��v��RXS�%J"���`7ě�r�/�������N��!�:.q:��z]�J�hH2B9���&E��D2�����Fn=�V6�\r���ո�8�YX:�v�z�쌂��n|�����~k�v��\����H�B�~̧���SU�q�?��/�L%��%/��x
#{lKӎYkƜi�����ɵ�2Vs�K��f\nܢ��2-�W�kz�;���-[I�́heI>��*T4�r�$8p�����Ĝ^������-��Z]�����eΦ!��O�Ρ��h���F�������n�X���:�Et�t��A�	$�➀����я����rcW��s�\���)F�����N�n�ߌ�\V/�?j�/4�2��z%�6 �[-����Ξ�+�@;%ek��á��F�����h��l�&M��.��$)�.Ǜ\��ͥm%v�|t%�Ӹpi1@)�,l�U#��̈O��>c�i_8Sz կ-!,2"�KԞ��h�� c�I9�I���ip|Y��bO��%SkP������R�a�q���i|��l�p�y�^�����3t�"��z^)e1�ˌ2��yqQjR@�f�b�\�/��-�g��M��$�����Z0�>��-��M��b��n�:�LA�˱3��+��Wv�8s��N�ETĴ��Jd�f���˾Iq�E%��*������e��M���N�U��fo��2���t��Kd�Q;�]c�E�ﬥh���N���Sh�K�~��8���pgh�_��c��X�?�N�pA�{����(1S��\B�J�ҙc�fPHs#���+ތ�s��"�6���l`�Vwx�BX��~��e�,(��t=�L�H�1:��T�S�t����C�j ~<��K�E ��FB��[EX5�̣a�`anp���eP�%���t�����oyp!. ��W^�Ӂ����9��k�
�1�(U^�H����~P�)��O�gK#�d#�oU|U���{�<�@]<��\�����l@[�Mi2�+Ўڪ�e�_%�
��ߩc��>?�rq��1&uPM���z%O��x~����	/!�X���&�(w;ʱ�WYo����. Ex��R�/x�KS%���&;��/��UhS����˴��Ŋ�]�*-�y �mF�96���77��жT�Ng1�-�n{��W#V����L[3ӊQ��9=;3k�0Acnv�J�]s���+�\f�f�LQ���K�N���5���c�M}_�I|��-�ȸ�X<?����7#~/��<�`h\u>�Cg��0,��#���|�_B��n��n\=���g��)5Q�ʯ�=YCl؝�Ί.��^��r6,km%�ޤ�g���c2P�W���F�E�u?D��g���P�-�AŨ�{��ť`�����șT���T��k��g��)�\� S\��T��}�Ъ�#ݓ
�bADt�u�
���H�oK�d-�|�	gi5��C����To�5)m��H�K��fPi��o�l��ڄ|�������0*����yeN��f��S�_F	��A�*�F�+ݕ����[���D9��#Q�vpsMu�sIg_��sTV?9�#}�W
��A��&?���9Һb�w�	�����	�We��.����Ow�i6��O�+���`� ��x9(�g
Ũ��/ͬĈloX8��a{{`���MD��#�p�;F3�$�*i#L�y�b ��̿���'"T!�l�D���T���������a�թ󸩀����Xv��k�;�\�c�@F��ҷ����	�C��P��~o�p^Rk�.�˳o��[[�T�&R�,]\A�S����X�{��[Nr�	x�cҊ,M��UR��a�ۍ/8���yJ���$P�W�;@�����\|8I�[8�KKͱ��>g����_2܁!K����Y*�X뱦7^b�
z>N+0�u5�%x�����uN�\}QЎ0��r����)^�o(ڟe��z�N��f"AA�EEnoE�:�f&l/�3��9moun7���ռ�Y�Զ���}|�x�|,�[�tB>aH�8a��˴.� Ub}�a#{�k�ӧ�D^�zk �U��"M*@�~�`���i
����ذ�p�9��MK���c<�SS"������+�u��6�3�Y��lQ�� ?��=�������y2@k��C�0܃.��x��8 dE^�/F�?R��m� C�NX�!vg&���aKQ�<Q��� ȣ�|yTS98��:����6?ʹ|�����Q}A��d6�m�o(���m��>{/�f��*d���􇡙��J�J�ꅹӎd>��Bt����O00֌sG ��GbS,��tQnC���B��S ���i�N~9�����zA6�9a�T��V�P�`C#��L,7��EǺ�/G��|3^�W��M K����}t�I����gm��v��.��G{��qQ��	F�%��|:��p,�6�� �37��̡U�aB�J�&+���4�>���;ûD>�5}������ ������'sͳ���3�����o�Y�܁,H��ny��(��nL؝jޙ7�}��u�@õ��^��oI��:�
6��"KA�֗�T��
��v��j������i����k�6�9мr�i�Z ?�����bPK@p�����7'�"��o�r�)X>`i񼅋>�F�C�~cJ.��0^�s�&��g��?�����Ii��Y1��BB��y������`��5����#��|]��e�4�T�	C�V��� �?��@���32��M�[�w�����#z��m.⼷�J9EuO���&�]�ۋ\q���	���K�5�:Ɓwa��3ҟD���D�U��TW�ZY�4�ER��l��;�//�aԅ�}�Н�G�q
0۹.5rݭl�y8:�o���8��s$�UcĊ��z���?�|#M�&�j 5�Lh[qG�Z��㸍���_ұSr�X�Y�V�ۦUs	o�'��.S)��₃$�<z͛��ƨ#�����/C�ȓy�T�λ }�`^!k��k�`0߅��Á�-K�Ju����pn�c#�@:�l�q�h�2�B�X�Td4����?ܮZeͭ���ft�����d�������AB{�����*���(�������e|OP���b�E~#J'�-��7*֧[��$�א,I���G���&��������n!Q��0Cx�'[-�5�`:�t-(��8�H�����u��,��U�ܷ#V�[�$�Q.3�1���3�������I���|���d�a�נ����3����&�
s}�0H��0��=��!0�����r���#���KWA������3�j��d*�<g�D:�)o�7r���J`4�a����/qV���ʚ���%���G��z�}�/�p�_�f�υro�Ff���ʂ�!�}��-f�7�<�������;�$���=b�
�$L��t���X{��t�̂��ed�{J��^d��>���r~��b�)2
g����N�G4�2�aa~'�E�)e��d01�(�2.�lGA���ٯ~��O^z� ?F���2[,:��4�&��ah��T��B�F?6����	���5��Jc��ҹ�ܱ����89V�4�=uG(���JNV�H� ���S�@u����H�=�gʼp�^"��K�̮���C�W]�Z�$�`0��גU��a��z�	<N����DH5��0}/��K("�o�k�`��R�	�?�EBl=����7��Ɏmn~�(6͝��X� ~j����v(�X���w@���o�V���,aEVj�4u��X�ּ@����f�Yw�����{z��$Q�:}�=����9��n<�<�	���yJ����q�LP�қ2.o�v06܆��a�B��\�4i��@n݈D��u�(H�������!<PRuc�@7��R��0|�8-�˘?��:<[m�����L�?r�?ue��#��'�F���ˈ��u��uɢ".0��m�^�N|5���$�ӿ��Ce�X�Ni��9׀��]���1�yO�IL�������Dslᰍ9�;�!_C�sUD���P�dO�)�9�,nXH0����6='��/g�f�G��Bg���|��JuӼ���`7�۴��Ti�;�l٦�v��m�(��р�х��W6;����؊�L������ω�@�-����1c}\�]a���t��F4T4a�|Ƹ�X18s���l���M����Y��-�S}�A���?��0� o��q^Ι�����$��A�1S���SӇ��B��`�3��+^�OG_��S���:Dvo�1��[u1��Q�pr�FFM\�6�צ����dr���\�&�~����zZo >@�GF¼��]��-�!�^a(Kg���TD��4�V*��ٙc��5�,js|-Ci�U�bQ=<��#9yfأ������[\�0)@4�A���x2Y���h������~)��S�ڄk]�\J$���a�#ډr��uĉ�;E'5�淚;���^5�>e��[���=��n	�c�p���۝!A�F�Ӑ��7���[q'�S���a6M���#�/ЧTK���~�S�<�΃�&5"�J���1�`�"
i*���� �*x��Y�6]��ҳ�e����X�ᙸ�;����4Ͽ\�2����2.-�ߩ>��/Yq�u��*{Q����`)+��/�[�z�Ɍ�ϰk��D�.Xv��� =K�G?�h+&2�����<����uxx�k'!=����������.5
�WA�)���Z=�+�V���~[���2� 򯴆�leĝ��Uڑ�ĎR?����+�&n@0�Rm��o#.s���F�������.��W� �"�缋�(e�Y�V� 7ɲ��Ǒ���l
JO��o���P����-4J�éW����y�=\"�v�F�[�E���m��G_:���Tbg���Qr��1$�O�S"iJ�9Lh� 6��E��!��Ȗ8p�+�M�;Ԓ��r�����{�����t���AL�'�茀��5q	�
�ؗO�]@�Y��\�"�	?/�VED_x�1<�":nѰ��t�+H;R���7��fc����� �Lζ�M�9]s����R3C(�3����F=�+	0&���Ğ��t�+`��ގ�6]@��*j�8�� N��]�mԐ��)�v�&�.;�T.��X�����	��-ZZ�����;�C>�����up��i�8Q�H�*C�)��J�f���u��o�w:ݭ�7���R�j���5�)�C�Ռ,U���Q�y��+_
����H��3
1u�y}:�������]مJE�g��՞V�r��~���y�X�`�Ԗz�S��0Oy�эO�L�e��
k|L��E�����[`�W.YP��Y
=ő��C�D��%����:���m-Ԉ��3�o�(!� S/�M�[D7J�~����fϧb��7�����:
���`x�1ٰKCa�6��9�Nӿ �-3Ѭl�_���?�F:A��n��	9��IH��q*"���z�9,���6�8�H����V�+�v���O֔��9�P�B���a8�Y�`�7�ب-R�4v�P5S��mh�T9�pi	�Z_�n��˙��s�n��@�����.k���w��E�@��uI��oG��0�gLͬ5f|�s���߻�NZ�1Ul ���QdL�I��ĝ�(�u0��/����7�W>�OV��06�5B:�H� ���ۃ�LV�y4�b���	l�N��<u�Jk��&+�sJEo"!QCMi�A2~C����@��Z\_%���C��8���AU�l ;m�H�Q5�<硌`��Ep�L��y�RƵx�D�نGJ�,�ݼ/S<`F����*8g��ڡ��jh��F�n�-���2CM^��Kǿ -��@��Rf6۾'����o�(?��H��wUI=�c�4��y�v��0��j��U�~��k�\�앗��oU��9�v�m���j����M��c���bLn��<`X����JY*`����߮o��+j͢�!��Z�K�}g��>����*�h���L�dX��ʍ�
q���%�'�4_�ʉ����vmz�-��ֵ�P�B
�����4Q�W���sAQk��p�.�iise8��h��Sz��7$����3%����['��l6��9jG��y�wt d����Cn���̳ϭ�:���]���A���;ʎy�����_�F���;d����;.K�	��_��g=�WJ��Y������]�/��������d�sn�$=�Q�'Pe��q�"�˿����J	�����F~f=�b~:7�Y�Psp�Ç>��Kָ�������p@5&�u,g�����Vץ� )���]�Ɛ�xO��}6NLa{���J8
�otr� /vA��wG�W}��{����d��`s����l�9K5�%5U��(?��ub���/ͅ�E�3W���ѵ���``�^*�7��_��$]'*�?2���<�s�eBP��I#�I���)�r��oj�éHd�ݠ֋�2nUߕ���i�|C�Pm�b<E=L��H�g8�u!u�6�`Y!=��z�l���`ģ��؈׃~//��/��d�[t�Ԕ+o; 0�7�&"��P\+�Z���?���0C�{DJ�5�w��=N'�`+������0����W�/�Ĝk���i�)���!����r�P�Mq�`?u@L�@��*�7��Ü=F�E�����A�s�)þ�or��YW$��3��9�Oc�����]��3�Y�)�i�r�*a뢱+�*���W19�
`�AA�+]v8m��_�J��I���!�_�9i�3B;��Ѕ�oc�
 ���e�?�Ś#^Ӯ�;�P��L:��],��k�F�4�82�ϙG��P����NC��T|�4{��1�3	<�64�b7`߳8e�;(�MQqeL�Q��`P#L���C�ڝw�̿f=�-icP���ǚyc�GW�uߐJJ�Թ���@)�ઝz�iI�i����9h5��x�M��a�����7�^�|��W` m�|�0�B�$��<�\HMX�Jzd,2�r��*x:~l��/UP�����C���l����j9���燐��*k4%տS���#_H�'�fU���w�͇ڞe� �/��L�R�o�57��~k������f��I���UHۿ���,�v업)��nu�ɰM� }N��0��U(�����j��\��6��"��z��T����[
b��v�4R�ŒήzdJLIQ�Yd=�*yr �k0Z����F
��lԻ5���C��vct���	u4��˝E��@�M_�ީ�>�b��3�0P4���
���Y��	����N�up�w����d��:�U�5�m���ѯ�u�ZՎ1�}��so���(:�z��u���!o$ $w;@�٦Z�M	�ė1:�������j[��[7���@��U�͚R�|K������fNz�ڤ�e�}{ ������JL��Φ�6,B��D۶�����c�S����|}��D�������jÝ&���h~�wÔ�vb�DQ���+ְ�c!�=��; ����-�������*�
!/)����V�2��mdCD	�2Y�Ur����rԥ���p���3A����TJ`�p�O�B�ay$Z�a����و����-dp����uK)]ǝ�-Ng�ߥʺ\k�d�ޢ<���-p����K�~25͍��L��E� M�����"�.y;-�-�^���h�>ҡT�6�-S�"%#��2I�A�S�8c�8$I�k�NSZDr���8���
����ax7���M:�H�`&�GH5i�V2�Z�Y�($��:��-^��e�����3�"t*r���H�	;HG������>�[��z�:�ux��"'���C�R�ѩ��������r,��~*P͢pZ�6&x�W��1���yh^ �&y!�'��h������$��d7@1�!q<yZn����,2v��'(����)�Q�Ŧ���uH3&��CѠ��R�^�E�f�Sp�I[6/"�<��~��i����[��ϞnN��ۅr���*�nBԌ��	�z�iKARC侼�d�z�{�����z���r�W]b�e��'�A\��%��SS���
CT6���x��M�y#&ZdI�ӆ��fz���Y��Q�G@����R$��Gpp,��89����,��j�x��I���Y���/*�읩H�j�9zgX�B~8�����F�2�����W	��13$�@S��^ЍSL�h�S^p��Y̅��.~LiN዆?
J^��F}2p^���s/E;,�jFm4�D>�85�?c�;��?bU��zG�n�(�^���W}Z�ͫ��=�T|��ktG�u�����$|¥X��'2E���o����~�IK��Љǉ��������Q��cj5�GRFݻ�A�3]�d���P�o�s���͕����:�	?�F��E��Y7����LH
��@���[�9gNL���4ߢ���)�b��w��I\�!N\��r�j��˰QJpz�m��a}�JO����ZK�+A���8�d�K��5#��зq�N��}��T�T��Z�#;������qQ��
<�{6Ϝ[��V�B/��MF�A�@r�)���G�˓��iK�,�7����$��ĸ�ld5hV�G&��;���l|��W�+��b(ձ/�f��ζ�ioŪ�+�A�{[����	��#4�ͽ���ȱeDi���U��W6�W�v�ݞ�/��������{'�Jaʄ�3LnK6:�("�m!�R�W������WH%.�&\G��FǍћ5X�zp��o�����V�Z �u�8���-�v�I���'�ϞN�M�h�st�ll�n^c��?�WS�7���Bg���_�Gz��Y�@�d������8%�[�^��7@Ӣ`eY��%�ZE�腿�
{�wYs��uu��h��
�}�$�PC@1}3�=t�6��Z��6с�sl����}����Q�Ju-�s�zUwGۂȉ�`9�b�ۜ��o\� �����T�4�F��sL
��X�G1��N0X���C`�B2�5HO���	�9�0��I���z���l��12��*Y�G��tR~9U�! xZ��b�G��u��A�b�������6��jHh\������h��G[Hļ��[��Xw,֙}
?q��\d�c0}��Դ>L�p"�%��J�F�&��-�����I�y���*q�֍��1G+@��- P�˨�Ƅ�ΈPM��֫�B�)��<�_�����+)�|ȶ*�(7
��A�ƟTTeH���\q��KaϠ_N�K�����K��".�p�T{�K_�Q?8������׏�8 aR�YE%�����ĆiNGO|�y0�m��}�=+�a������a����8V���3��������u{�,Z,h�KMGt� ��;4�նo\H���D���",��z �.�"By����$(�]4�L��yZ	G�9*�V�=ߢ"�������R��S�r���E��^� K����S�ѝ��j���	�Աw�.�F�!��L�;�� ��|�%�,;[pՕK�X܊�\����'�y ��bBw4)�M��c�݆�qV��qCϋ�����ӐKz�S+0Sӄ�w��8�	�	�RK�w����|f?���;�����ͼ�֊�s�_�$8ƛw�����q��"m��ɂ�b�E���j�K�Z��D׶	]��[�J)� 2