-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
xTFfXah2mtrWQf21+hRZXZb3KstGCQ0OiUhH9cT0zqSfcVozn4mMeVKXxb5afvS9aFF46m9k7Ilz
yFT+iw+7oraIwvZTGiKqPnufXXOLAhuD4GUFXnTmrkpI1G9Jyg4gPuQyPeIKG1BdwtqBVwifrfBC
UkPQvqDIj+45ZrUY+WM1NvzhHDrQeVoegWyoUGzgJT3tFUDixzh9DD9XmdgNNhGC6x//2CkA+LRv
ywBPb6IcB6A/EgIkpAUZ3wj3CjVFR4KGGLmnlzo+WN/HvDky+foL5lPBhcMTFE7KZu3FtRR5stPN
V4XyWsNcFhgNJ3tGLvYAGc4EXM0auHX2A+NYSg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 21264)
`protect data_block
Y+sIwa9r0tQsuJa4TRiQuMMZkDy4saw4VMZ0S9ZZKl0g5eiVzJ+nNhIl5+BKMIp+MhJ5dm522/jZ
H/+SOSDqc4iemupdldeH0RKedt6d8Az9Xq33lGCwJItcGgP3wsmsCKUcLykk7Krr0XEKSYxZKmHM
Kit5HtR3HkENOpES8rOT0tgf7mVm0sgJxiylQzi90E70cqRFxDV4giDUjcoj7L4a8dnwKsYMD9Kb
/0mcKbEidFiKGzE3zQ+O0sMGKlc2D/v7BiM25PryIumw5KtgAarSJEhVzrOqWv7W5MnoIWEzzQ0g
eos8F/5tA+WVNo2VxAYL9VvkWcpFgk8heURJbREnp7EW+7iRYEF4Su4pBCnlpG7xzfnlQoiCiJ5i
fi3F44rTQUhBkpbqH5Tdn77DDqU7ItV6BUD3j2ZxNsef7y+l3BAppeXnRu5ATqtWf3VICkwBGlcX
/WDh9VYmPTwtVDOf6o+XSwrCUFYWP9Z5KXzC0NCexyS8x3+fg39jCpCWvVtA+E/F5KXN38Nb2VDA
QRmIPh8OY+VvrKeCwu7OQh+Ox6cb4qBYssn8c0QoRViS0dgDx92sl3FxAFaGrsa4gNPv6cb7hdIY
2L5KHwytmQrA+SnelvGPivzou7EJHxeNpLrqVAhp2+OHiuw9paAXSJM40+D+0O7DdSLVChPN0ryd
fz7QZbNBzixf6vk0p4N8Rc3r96cXMMFPsDfQMIjt3JT2RrRVhKM5CL5eVEWpnWTCmgNzvyb9Z3TD
xNUGXqEFWPg79euCxKofSq4tnF0qP0Dleb4W5oUhI8wHohmM807gfprd2HphKoqYJ28E4MmGosDD
xoz2fBPZGGjSE87nd4SGO7DVfhHkvZh+XnV9OY2zUOb5VEZEgVNncdxsDrqcbh+E8xbeEAJ7ByvF
Hnwj0u5jhi4jdURbWsitV3vICixJCoGCsuedJZHSY6jWmXUFo9MG4gKyXKqsIsx7azR3jWX7Q1Uw
/rRcYPxk3Qy7+h8+X+OnYcy+aXHW4cmvc1dyFFo11X5kKLzlPz0XYaaceM9S6JWLYkBCta7XgfCu
Z9AlCPQR2b5gjPwZ3kvQgWfjXswkd23Ko2vEcOxOrTkkE0pAbDDqVflR13iP/mUW2XsRWPgsviKa
dCU70W+Jh6WLgkbS2M3H953vO5UD6axFkW2xVNjiIpeszmvW5GqKGD1M1WQqD/w9iXttZYlWBMK4
F8XNUJzr29L/8Of8ICcuUZlt+fK2HkwbIN+aUhCDfBn5VWg3O7PJ1qz6FkxGHnhiWe0LN3XbB9SD
QXc/vFl7HbfFb1SesaiFdGz3vBkMy1TEHpte+kygY0RW+9seP7oCjbigNTii7iuvi5VFfkpvT/3u
qOexYkkyypc1ut5ENnGhul1iUHYluODB626Su01/PEeUOXE6Yk0UdFmH+Lgk8NxDwFk/54WILfY1
wqW/JgcUvWGwysZlxzaNyGk+B4JC5HewL+L8ZytHvR6xpq7NlHpEMcy31NmW0F0T6f7tP2e7BrZi
FNFZC5thEV4HdicFfwb5jKf3tNoozTFaDnRVx7OIFSOP9/aq3fmu2TGruKLnGvoGfLHEXxT3XWvY
Was0atoq/+S084arzJTGttp6LW3Gh0csUC9nkocbkjEM9MOlLYMdRT0ypb7qJmMgwkVbmzLSG9wd
KbTqbok/T/n/b9avLcFbxeYCjXD+L6lXu7laHkFopwkShQmpky02dgfh65pZoR/y0wZRYPA7ODcN
dvftZh/UGhwlU7LAU5gdK4JDgdhKlnFBF3IWY7F+hoEd/Unk3wqa9OHpL1SnUUzEc7FUW2OAAuxw
it4cEfFKmeeZfXLrG/90rBpwj4hXGtp7wUe5DVS/MU3M9vdZ72AusMogfA9JKfDfP/dsvH3s3D/i
MtUW+KXM3+qkUZg3fqJ61p+odPU/JZXrNfegQsBQRul2Lkz1Y55Nyn+ajKXKWyTx9UG2lBSqWFqh
qFXJzRx4RkD/8yN+h81gQ2hKoJeh/KtvXmZR0p786ybllGLSXuwWhF/ZjDCn5T4NnJhV6Zn4+S9S
W0cCeTHGFp4BeHtQnV3W4w22eLsNd/249G5sf/64vDd5oyQa46AhfBRLXebvoSYPZXgAT1Vji9TI
KQlQzhW+gQ43kivorysRRs9qXT0I8bbarM0SmTbxyk4fM8sfW8DC+qI4l3nFwiVj7WVWC63beQQB
EVcRndpNq40GeiN/ml+QuA5fgftFWTrn3BxkXE1vFsUx8JPARO8OrW+zCcO2t6AjT92OQ4dkqsNe
MEMzbU2Oo4vxGPtR5WTp48/SuNxY01/6WuvqUwDg/A0bbNWsuSRUGHySttXp3/MzXFmqCVR4Zc5b
j7zd3/JYftLBmtI+QlsSEy57Yq09zue+qsJ5LmFmajRQfIOAazw2ZfzKkl2TxvQIB37Ju5+uJeNi
2bmP8dzuPafQe4oJR48NV2xbbMJ0gvHhyNsv9rqvv9IqGEBJrOLuSfhawMGx60fObWaq1jSI/EEi
474wx33NJnPnFP2EX+OlV4Mu1gE/aYN08LJFnu05D40ilF+BAckEpflWRRJ2rs9yVVMCDGo8vhr7
oEoMrdEgBxxq8vkKEUrlZ/8tgLuRu1K2Mb+apmNlPuD5oSM7ovle3AJfNRfTzDxg4tqL3eR9i73c
2BTAvENmvYLeXmeSgSuPijRdQOarX6NkfhxYbdKGTltlLlBnEuMc8WrugKohvJSr9jVJzHxT3Ov4
GXbFDwwG5lblnuKwkaklaKohGhoQcK8rfuCBkneuDECCDcjEweCuWXC6pUTXLyvTE+ju/y96Poan
Sq19PNt/xaEai4znnKYxv9eUOleafA0p1YNJ7OngiRDq2AO2sO5Gmk0IU7Rm7InMElYYqTHaPw1r
a0LvzoMiWWIvWXiMcf/KDmX2ySZxFTQqxnC8ahg7vFFTUqA3UqrPQeoNNKtDyJlOzNdwg0TkN7y8
NV6nv+S30sbUxFBygO13o4xd4z5d9a5qLrHRcUCnICy99g8H3uIuMmY2T2IBOHdkmBrzwrp5jvks
tAOah4VbqbcBnHVTAr6fDO4J7LaQt+nyiIkh72o/9oY7MFr8Vqc2K8g0v2KhB0+1eD5awuEokEbA
5uoIKeDmekiDXMnJLPgnwdh+Ew0YDuLgjaCkgRsgoyTjhn951KJTjXw2QyFSQc+dz2KoxuwkhnPS
0qBTsprGNYpavow4Z3l8JHwS2QBuSTSSEWeQRVCAyzJZTL7Zj7atKv7PChQJG9nPukqOzP/0RqyS
ynsjgiqkntrOvGdxbkKYs0WxHJ/v4so8Y9PPA9JUsjgpgQ88Kw70X+014oi6FmD63YnpRLO7zA3C
jbPOCKHR+VmkbyT5imPN57LRqTQedTERsVWZHXF37ZkbZwBR6zqwJV6BiwHZP9sj0VjLF7ICgRxO
IXLjmkRheShRcAu/HaNtXegXQx2ebNflOCL+HrajNx/bhX6g/jJRDSpuTVHSI68RLfeqcACpIz+L
S3M5t2NsdgVoyol0FoFJ0qVTLRwTMXdA4GrGpvl4lPTgFIC6qxOYfsO1Qyi7QopUKMRlt3hxka02
Lj61KsD4P/QLKsYG0LbbqJEtBWF7DYyRnae39P/Cs5ByD5U92gRg6Yu0NAdtLdGxZ3wzxAPLkr/a
8EEawAzJZ90nbXhDe+I1LygmfoHPXj1FSGufIN5FsFCAPY0ltF4sl+A8HF42ZRMy4Q7mLiXpBFgy
5+v3RBRrZq28QOSRs3k3gpdkGRCQFkiaZniF7PMTCXwM+Fhx9HgGPe4dmCeysZUch6d+Ba9j9Q5G
t5snvmNY9zqoPAtV/FhmjCN1SfTr2+LpR5yUp6ievU5A0Ennb8HT8pcbjDrv3Tt8jpZc9D5FdbIl
YPSVcK+Cekk4z2ZaIf7nsLlYF6+PaUARx8ezMhEtDa0fuG+h0GgdzvSNzHracsFij3oLmpSL2xP3
3RJOVlE03NLxCAhrtgpyoUgSoZxn9PngjdnPNIxh3zRZ3mzC3m0nF9jsvLa4psAfsIVd7WkMfwNK
8ktTMzCrPGtMOWoOcEacO3alSQP0P75hksInojaS4zmvfU8HEfshPyrRCF4WB0eYjzxKrFu8Xu3U
aAJY8y2cbRvyVA7LMJLUabGdBbhmJs4H7NwJVw415NScpIHN+4ZpSZy8S4tEkthJLXkmZqsxyqOF
zszpGkVu1W9Xx14wXXmbg3QG+Vvm57lliF39EPqUVze1FZMJ/Ck2OB9RPhFC6OrfEPisDEHEcfIM
AppNs9PZgHmLy+xSeszpoW6VllkOlkI6nKSwA6GZ6mdLDs7woDuRE3TVzExYrPZkYr7lU4OVazXn
6wqv5E95LNu1S4PF66rDo3Ko7FyekmorQ/T6segxcnR0FynE/ETASCUBTOF/5SwRhPKE4831r7hA
ExQ1cnoWg2qZPk51fFkDalfjj4uuAYFk5N1bt5wlRyQqxx/b6yGmZsgP9ih97K0BgKy7KndBJvfl
NnLJmmykX6mso0I5eAt+2VkvfgxgJ0ZvhCVYwG2GtPNUtlgPon0JKCRWNT9D6xdbSQUdtprziN01
LJQaOrUombfJfO3mClbebgLEUgJQJzJsg5FzfufzkCqkWbWjMUoWgTnTf4Isrkd2gQ+GNgFmqAvB
3d47rkoLp9hRNrR3236/v/s67RgNdCJla4OnS+UI5tRR2mS7nXWwC2+PmPJdZBNFSWJB1NfSaLr4
j3ST+MkI48GGqrEA3YxFxcefrxWtk/RtQXBoeqPY5Y8f4IKdnHsIQqdR2KjFZ6e1HI5X4CnKXrGq
E53gqLLDw6z6VF5Y4lh0ySPvlbAnqx5f8uO2TEHrfuV4GUeje8CbgxsmIp1k+dWyJV9uGxTETXdy
pOccz61KMtaEvNAjRCUPibVyIJL1omTBeyouz1GlkA7XXyojkhs5N1KnNFa/9/2kVuMTRIgREdpi
aBo67HJXB79VkCHON/BrC3MRH0BnChO/LbgWtm8o11efAIyYsTRoEo/Doe7Ab+maU6A/AtsigpLm
iBWP9jPclWuOeciubYl+ZSwzu81IvfWVB6VlSFY+hQndfG4CKlhzsEMhfnk/H/PtIfdA5n2jyej9
IbOCE1axNFqZZvPFQxdmekdOojabfgdllrEES8RbKz5L/fE+HrQ39OhI831gy7r6hEuB5eeli8nM
s0yXBmZJhrsP1YEm6Nemah/41jAZT49qLcJug2YdDSGuiF+IABJ2pfIx8kDzNKUOI/WXooaQM7iG
M9plNjzmYZCr3DZDhQD1QTLyxjZIldAiOpn71NnLySMZMxzm8EatvTWnd0fHMW2R+tnkXIiFHypj
FmW8UxSjSGlJgymPsvuu/AeJRa9LfQWeCBQEnUML+gdrzlu83ZqE7rn/npRSkE1GVpvA5bz4BP10
HycraQfuCigsML1q2gdo01Jvx0YmucvNYeqDFE4YZiXnolgCvpp7Pg20EwyFJlqF5RyhW7gVSSx5
Fz94M/yghfheQLOpe9cZhBwOIUAjURMPGv3N5QlbYnJe8qKDPRNfFleUCOqVGgk+VG1OrBmj4Cmz
iiRVkav9ZmDPMOVJIYjd44uq3+/Ja/aJGLipdFlQLXF/64ajek9iMsa4gbdULGQaev7aRLiLfYkb
bPfqvJSl8nx+jCH6LIY2YBuA8JoNQjnrxfaJXzCdMXLBdlg253Oh0lEm7PmDO5jJjJ5LcJ750cyf
LvmRO5YZOsnMWL5adDwyMOW0yfQYeVShzI3gj0T1tjd9ZpLt1A8CUUvI8NrRCmbo4GgN0PC/W9Uc
PyQ8thJ/6XpKQIpTrlokM47LZMeZap/NrAR3W5tk6GlZJW5I08vm4oV5SMqZuLeOp8VdHu+7BTNd
yKBMzJTvANjApBbGmLx02Uexv46Yd5FTMBhyCp+deYaPzkvwRdNhnHPivKnUW13BuSuQTkIpDQdh
0zslrrqpk7PtRnbD6qaOcQ35OmXbxEkm/gIuws0L+G9vYbcMS2xrLEwr9ARnGjFq4GGswvoSinKI
NgwtofcovNc+asLh6r+cqhp1o1oKHCq8qR4enGLj0kAm1zY7DVTWKoZ+rc1BNE7B7/Rw/7zkWuxG
tCmS18FaE//FGSpRIIK8AZL76KrncAHuKCnEcbMKK0lY93OjVVu9HeJaVPKWwRDMezT5uEoLwGjg
+5PrB6R0K6aJJH/07v7dkBiB0YRZSvDc2JvzN90mtzYkTXziOSkZ0bsKzRSiwj3OFqvAZrepcdsb
T+Qf0O/vPFMg0bAlWf6ZhDUeXH6chXbA+8qowpCYTFuWypa/9FHn28PWEu7L/IPfEsSIozrrXVWL
EsneJJsABm/g0CNTBGKhc9BdowlhTZ7hSKHWKKJEuOOozeeiy8NzGiS2cVb2/RKOH/b9h22A7jiC
41gIw980xvm4+fp2PSs6SM+HLQD5fPeUjhqQ5l9xz/XawAz1/JFLJAeR5vXg7Y1cSjunKWmwKusO
ruD2I7IZd9pb5ThCtjnbZLIecqCxfHBnJGn6IqmawOmIV9pXw2weglPEwm1ksj2K/1Pu9LBXzG9N
tiQP3WLJwBnbBlxqa/3kbNNg97njKNWyOKwHbHXqp3E9AGDSPUsD757ieL9ghhS5WUDXyIuXYiLO
daPUSP4pzHOl+8+NAOSSJiOvI0CRCnumEoirFwyVawO0JNPe7DTfe0bQ+Zir4J3pWOtqv/aAKNFh
LxQ04EYK4lb5F8uoZGoQSyfy1zg3fy6eXMVTspfcXCC07unHM2SDG14OIv/aoUc6N7SP+hfYbemc
MrSV1WQ8fzpt9kSBbBH86p1smrSqoOV7rZDx1yJNO/Y76BS+OPzTw92tRLF+W8oAbj5/131qusnn
IEsUoKIXV+RhCKPauH9UH28Y6A+SMXIHdmOLYJehu6j1JHeDHRGec3SQ219zJhx0+X0jPVXfINxp
AiBWA4b6qVgKi+3hL+Hs/Gvl/CsoF8adsu43SoF5bhl/cIjbCdJYAS2ayvqavxBJoiFZA9Uatgow
ekUrNmziAGNXtWC9YLy2T6AU+56rxdiB0cyuFiPkGvc127UdodqQCQ4oHUtl9KMRUGQUel44DV9W
NGIw9bXXEyiRJOeKIEcjf4xoSMqYoxOuI/iL53roqgl/F+velii7PMaE5K1PfgS0A1QK1xORB1vd
zdA8mSt0kvi27y8TtUQ7eWTovpS6MB3wbzsy1INqGKDs0yykjQrYaoOLnuHMLdD6Y4hY6N+Ccsbt
dXF5q1B1fWHi04UU7CElaaJaT2lT+uI1NEcYqP4WyPf35vSL+6rEqd7UKXIeJ8iHQ1knaVyo4BaR
/pNVAMHTs5M8D3dzO2XLJf15nxN9cZLooqNgTh0xo40jXGd7GusISTYIthFyej4iiztqeTSKHc4k
wzNma4kIv+vtRvm//ti1fTaWeboYe0aH8z5x2H/KvlJizEetwN7/GwgSLo7lUcBBqHzveUHcjV3o
gdoVvtqn/DJnQCapxv15EQ+bnKown5OQ3WD/SUYcKGc/bhjG/YxMon/AOw5dZz5NDWY1BQq8ncdf
p+i/CKWH3wbNg39yyuGAINQ9gvROz9TT4EbHClZpo4jNeQLg9mM1bu7HBZTMlgkU2kY+yq8bGxhq
B1LYq6kVa2ox1h74MRrj+G48FoCXxp3u5Hx+GiY2JPn7GnNstcsacW6Se3Jlr7bvRBal4bV9mAgq
TnDZDbuwMqvnOooFFHEhBQZXKhZSbX61b97pLEtb7H1982QSdNoCLxdquS0WIYcMYqL9IAnb96qf
BgaL9FLsQi9om470qKILACheTKMsxfWeTe9dZg0V7OvbhXyLJNGIGIU7w8y1iTFb92pX9Ohvg8rw
WqLSxpvZsPg7urqu6cSAdoSd5JPPiMHNGdW/WRJBI2Z6h6e0bvIrEtbUCzVi1BHv4niwCmNkDr4T
YwT2JPkkHUd+5njLHdDOJMqbZeHssqcx2QEYAu7dBiRRvrrckVDH1sv0Nsi5hsx3xIvvb3Ln7SOU
bfILOpUINVqDcmh5XX6RQOwcJ58jvsWp30TTumVynmudH6OFVBHyeqMngaGXROaIA+PG0tjVl4PQ
PhIaBvkBs6OeuzZ+g3c6e8LuqEfEywsUOfzwiKuqhnCtwhN1YEEY7+JtrQe5WVRkf1E4E8FcaB5H
ZNjmo6NqIeVDgWcjyTPxW2JUOZis25XMNJqSPv/C14vsh/9w216LTkKIkAgP/bQBvl30OBfcxuhR
EAkFfxuASV8t6JnhegLfohPDvp0S6vFZc/wwh41EWHPs/Rf4dhYAjMBNyMjZ1aFlmsfHcOYYgqdz
4545ADYr6O9g9UQbeghZcNGDrpzBONiTG/qlUTBmBXCe75kI8Lm34zInL09LLlDe027MFvmm2NkY
ozIj58MuTzffK/xARSQEnkbaXinwORZKojXGzS6KE+gy6HWbsQdRBxTMW5vJKIc9PAIjdJBOmy1H
EpmZzOCwe2bvvl1xCUtm7bBrTWqCEj2UtnF+67bXLMoom2TjgdH8nmi7BbU/ZqHVD7OVSqbRm4IG
cALITy/GO4QYhOrZLA0uXcJuitkcKZMJT8n5lip5rsM7icy3hq4PcgxS9X1fMHUCPUrO/nl2JCsA
IDwYRcs2Rzuj1gJ2Bvf7JKHc+K84YjdBAg1H3mRRVPzLIv4Q3TTjdGhig3ezKOlVSPpJm0VWEE8n
YfcEIPCkRB7GCs7t/D+Q3bMQYv0zs808XVbcW3VYbk6IJjkzTVzslQs45mWqxqB6CO05Rvz7Be7L
A7+lB1Rn15TN+HFvX76y2rZ3tBXI/SnhMiwdCisp1CQxDYphcaX9S4cmIi3Lg32l6xkqgJOs4DAU
zTdwGwxKGHleGl3GFIhurdL7Rg4Izjj1eHYnFbpoW9EKX7fGeaoXHWhVAHUYUa1Vs7pKvKgmH4WL
Kr1V5GzHzSvFWfjzEo7h8CQbXIB5l2aorrOxIvUL4am5a+DOJwPKT3NYXdh61km6qrHnHoYSiHgy
f8VxHf238wXKNUFFYsbQPKO2qK4SfSSzJxIJqHKAHTqAt4e2JqcC1tjI6bZpLCvmpMvaeBFLsArm
nDB4Mt4EGmYJCdknYfaZR/c3hAB+qOZkHC+xS3PQXaqjfG42HxPehAacSbA9nIyJVXHayfsxgZmJ
LtBivlJr/jK8dPWzzNDo8d84DqLoESLCQ+qfWsL6d0sc4AHNq9l5F8ghKLCCLkuVoELFL2ampHq2
gjNXphqXdxmLJ0aOh2ay42VzYQXP2tUePbWuEiIHyR05Hcg+eLonGlQgbggN1KRWx524Gk77qIaV
QLnRkm0E8aU7uxFCabEkChCll29eUDyWv8Qa3Pjk2mmDwPhF51e2EgzctitHEY9VJOpD3EqDvE76
MWKaVRvhPqmvebY6Vus+El0m/QGRQqSkkeKz6rb8uMcKcmvzUH+6NAlgPjZ371H5Loj2Z6NFbVaD
E+NxmH4yga/UTO4sOf4cJXwQn+9jqOYqPAntSxT0YWgmTdy4aHpoxQMFAtyKYg2ZDrlj2A3RBrLl
c4moGGXkkyk7p6SvMQYLKSrq1cTwagsYy7EIZriyGuz/6mX5n1KQoZNmpdqmrXyk180PgIKG6ZT8
ef7BWh1YfnnzTUbBccvz+MouCpaOEwKxkxTp8qwQyojkCyJ8jfXtNhnlKWQwrQ2JJU1JS4pHxgdo
5JZ3wBlJo9sFakgYIsfjmlbT4TYtHxs3QxTNb40D3y8WLBznEV+xaVr4ptiwCaKmYe9waVJvMRNr
CyrQL7f83m+i6geylANcFxagizBHBRZ0wwmmchvY+jws4htyOOwl7oAMgCZzRqAZ623cs/eZ1/GC
sdoY+EnZ1kW5jKR7ZJ+ohkNdQVP3TDLvjEaVtQPvC0lvwD229jK7OP4VUmH5E00H7fIL+lwI4KL7
nQlHhGKKau4w2rijK0Y6s/W7z5/5+zYSk/V8YwWHj53rXSUuXVs2pmvpbYNOOvX9FsfD0FF631ve
BQz3/F1brGYy0c3Ev6+Zk5g2+cUa8mNwZlUHW1GSdc9wFbE/TRL5ZAQHh30siEfLE2BbIMDFn5OQ
2rtAVCYJRXE4ZrOaeqq8pqy2lWUILstcmibfE9rvK6QEtpu8UyTMNtOASyduUe5Gn2ag9zAozUja
Iz8Q4tvhSq1JK96VHwcniAmwSZbGVBc0aBuAvTS+G9sy8qxHOG0MoU9tZRpyDEps78/dOHVnjX4I
r5YmlP0xPv+TI+GqrtiAY7+h8gtDB2W3ElY4Hg/SbkR9MCYpxCMmopXSMmn9MwSK3fyhU0cUzHqr
cZsATrba7AuhHNaKGGoaDnO2esh+qdcgKk559ZMoBE2v4GCBiVEa2fxfXUs69ZaMndVKHzSkdcWH
hZBA9B9NFoB3n/rfVji5yNbfXbc8ER89ImAqHZDl9qneXKz5p1uWE91nl4LU++3qADkZnRnkYE/x
ifE8xp8B8fHiwcPCJywaywOpqPeFm7BN1CWZZDir26p+vf2OaESBx7xbRXC1EtM+hhsEEMVcOByK
5lbevxrwSsKX7OEgAHvjGkO/HFFLQnQA6Ew0m2Wd0PGuTKtFEcnq8/lV5gfv76gl+liS2dFUi/IY
aa+1BbqlNHqBUwNnfr6Q1sGNMccyfTZqja2kK5XUSGC/meeqqTKenm+sEO8zMFudhHc0EYMmn/hm
/rCsP1eLW1ZyA3Tu12zavJuM+RarRER9O2gznjH1IFKfl5LOBimp+TSDOD8JxVam+ANr2/RzCHn/
xfmPmRrh/HGopZiep13z4XrtpvcY8B7hGFQjHzVIrNDS9nP4gihjgn7/nBrNAABOsgwcnjtsG5jD
i6PAg7n6HjmOk9M3LsyD3SC03sYwm16gRfZ14Tc3Gs0it3E0sskDbw46bvZVkTtUk4hXIKS7+97A
QylV71lzEtiVcWRpfb+4xgr40hKUw5C19/XFGhGVUeXzFfKS+ZG6/AE3cx5phqkevPOb/xpNcXY2
cDjkagoVzDB+FUqSPoS2pn0bzscxn1S0coZu4DvC1llZ4ne4rL/91e1yNwi1WtOlTYC5yH2Plb61
ibkYOViBdZ6Cal8GJX/6GBkuMQylr8v2udFhw9bEM7QWzOADZfk0gKV/5ywSGUjs100e+U2lDJg+
xRGojmr6vku1HDD2p2hlLU/HwbTnaiDt9whro85j26pkgE3WvNV9cSJRZflr4STWDu+HurFyG/w/
O5FdO0CmFC4douvkMaEHVpgjGwzkU6ho2cVv8z9Z7kpzs6hEE/MRVEWnn+UHPtC4WgXZ6Am7i927
OJ4jqT9fCH43ME0OWsPUE/81LRJezCbwVkYimdY+qkIz/uUdHh6gTFw8Ki0/RBhd4F6kymurjPUC
XQPmAV+9sGfejRMzQ/Rqv7UunXV33REbO4Vithk+5W4GVsqPhCYua45yEjkTW+5t0ZX7X4liy2gv
Ba03G+8WLIyFD8B6+MZjoan5P0mYu4BnwJdC+rlhW+zGx+iEqLjo11NyR3woydADD8sdKHZkQgf+
mm9PQe++1eKNm+FjOTTVw61wVLby2ZI8Mq43FCWvNCOwRlQJ8HPbCJcUX2PZYg8IZvzLxdLArUmT
m2tEQV2vpjwr3G1bTi74ThtTLYOfBFX1GTBCKIVBb9/4/xNleyXLmaszxkB0dpFU05LrzOakhxHw
R0sNK5oWbyLOG7dvUDr2a6ZJ4Q4yEF8lnLP6kJKK++wSBLw8jJDLaRqEMZawZEDGQ/YeoVoqSek9
3MnUwho8ELGavjRWYi1s9B0HY3xZQfDAzV1QzeJDWHuNEn14YVlXqow+j9hYaSjhVFPkVlb1Ng0W
0vaCeO07Hw+b3IVhWxNouCB4qGflOrDXsSJmJrOwoIgsw9n+HwVX6YVKJBMVt0DETkub1KAxDAVD
x5MEVwySw2zQ3rpggRhQ+4lWpbv+1rilE1jw8d4XcE2NnGiSw2uMLSrgzn0C3q4vB6LF5zvKHqLl
k146nCzjqDr+Zlp3l0a3r+bbFYpzmRBDuPlR223E/Vvc79YLLv1tvB7YejBDv7q3AVsbhKmDMp1C
rEGTuEwY+QpHwPfLlPBpoAdFuJYEf0PSQ5qveSZEdf6qQXo8IZH28SJWyYdTXKHZKQ4UYO3MZgLA
BLndz1anGnJRL522OkG85LTvWG3TvsdGi7gOThpc0rgXZk+L1B6x4zaOmN7OhNro6gSeZ9euYg+B
MQ7ahR5QxytxbcIGGNXa6SOLKVaP8vWZxKANX0sJ3CX0qlnJt/hrKr8jAFsEynBdUkU/MrVN96/Q
kGxEQFch2n9Ggo278XzhJG68QmvzSQ9NpmOPDo+EuDVCLaxAOyi+GuUXiKKKRMT3ya4rJ+nOi9kv
BoIcU/cbTHaPAOiWdedO53JEJlHwVj7d0Up91vrfdausSo+cSgljDoOOOIN2OaKlH8nZZDO5zYb4
RN+BfcLDQV89cI9+UPCuXNxjMNAb5XsF/xwApb8Eul6CMkEtaHbvlpabftU1VBobQw9cmV1CQX0r
Bz8LFAW/lUqRJ98sccf8+82WFoYWM+BMyy/kq4RZ+uuMfjKIxx8bPBE47XMFS9FU05JTLRuWZkeN
FRFBfQLF/govOK3M0+eiyh+zurr2LO8Lo2urXf6Cn1WAzQsSUBrgVmnqZNjF8EH/7zE0RxYISgPx
czce3oCjgoU5COZfXkDCxbDZFCy3gm2Rh/ADevKLcebVVpeyXEinsAKoaGnZbHMGbDi3ddzBYRlY
ZljvQrKYXKRwFY9+mMzzdfMReLfYvp8sX41CXMdx+SiIxPl4AuusAOuZRn/KKfrZ+mGZKJ2fDtIL
loxrHO9RwJQKvkPHKTizD9QIamEfVsbnhpsS+qTTW0Sk6KCwkawmPzmBPNnsaJbxVQB9DvMlNCuc
sPnsiTmp7l+CfwYCnQ68onFVvBlAAcVvdNpMLY43huSwLLIJbS+RfArsSP0mi2BRQAos/V71/A1J
hB0bcdvWLn0QoPzmhYinA4/fxfDIBIxgu1GuKjXvTxznGQ2+rZytb7mwV+2dXv56GDbTc/xFTujK
AwtmRpxfFHRSmKbq9ImV5Qqo2JS+oEpLt/lNd8k6VbhN86T4yS8k3Y4ub1r+23WACFC0PxRDGAfc
Ubra535yJFJg5FuUaXy7LMo5mLBCEd0OhP5qdLXgQTQYcQFyFrsfigOewj5b4w3HVPf9KJ57vsmm
qvlkmKqsuj48O+jyVr13y8x9q4JWB6qwgCD7Jt9vNr8n/5b3G90Su4AofGs6parZoPVeHv6m3DR7
QQQLJ2iX0cS2+r3cBs+LcgayYR05aG23l1TC47lz/ZzVJ/vxfhDRGyBmbNoj98i7fwtAO5H00qD/
prlFislUtwyqN3lSJmSR2vIdyQ1a1KcMGztk6HequOOg08043BNB/qa8t/EZCRTHTlgtdnCsL3V2
5j1ZHyfQQHcLXav/mWRrW2s4rO0eANCrTmnlcTIhVFXJmAgmXmrlXFy1+awOOrp5zZNaPUXepSdJ
b7Wv5DYisbwW7rw7iM1PXMnakRvQl9rs5bbtj4boGRA9K507vgWrfc6CiYYBOFIQCTy0CNyxEmQY
g6G4GBGYJtbahgFVvjtAz/p0hT0rizd+2Q916tTO8h8VTfzxShE0fse/CdZqj4XCkhtvuXDR0uMK
Xg5xvkyxvo3iQIEJq59B4gySGyNPuuGkmuOJpNa0hOb3CN+kKwpDDVLkGzv9tST0+9BdtNA+OiQ9
vTuGh502Fx7qBddwOSArSXnCeNAI/jwGmMT6FhJHcl22qfBVubEvWnv6ovjMooSFKkOm/BFYVnCj
KeikZI21yc+Kp5tDDvwppKhbx3dpnxrpbGlYHmPF4+u3u5KaNwHbmKdALz+QXgottCv7di3fkC6d
Pyp+3PnH9M+cnC1kJ2LB9Nl0TEOW4tAF2HvmQPhOKl4S3DUXZt1fhQfTYQE1WTAj72hem88cfUpu
K7B/8i8wxXFp5v3mmnBTPB+feChQLo72j5gYN5Qre3ra1ERSm1SF162UMwXJnHfxXUIzEQt6DOJU
topCq3xs9lXxD9aRBIoe30/nUpT/JHh7Wk3W6dYPLn9CvtrX/6UKy1Ri0TW4rsglrHl3SCDQy2qX
hd3eBf0kPk6MI7nuHchFWXCB4ZVrdrLHcnpjdxDMmS6AWe+8tD7i+muJdQYLdvBFZOzCy9IzjcSP
nqwW+zNNWxsC9t2PiJHrjg/ykWp9ZKPer09MP2Hum8zWSmIBMXgA47hxkvoEH10V06eoC1ePkfYo
dbDwgV5W68qlD5xXfzkm9wm+UekgIMKlou0/96aqzckEZA7w56omgqm1nUFL4+09yjSj1LHI6XHI
N0Il8Y2qxI8wcsdqC7IuXcnCiD3aVav26HZfQGsXTZaHVaflRo5R4KfdGTJkbRgxd16WUQtcxET0
/cZTIhKI08+g+s0xmRBL3JlLdJ4x0RUe49NPo8W7KAy+1vxrZXzgGnd6BC2BswArNXjdWT1nYAeX
N3Q6aiRTLzrr2r6GWdkhhcE00sr/D3/ZLzM9P9dl+gfL4X8mH1dsuPI0elgMT13vc+5gYLyJ/cRz
kUdbxci4PB4ZC0S0rn8aoSXOSE6u5qMyRNweuEeKSp/cCz5NKtJkOvl2+hCy7AxXc2uNMdio5k8L
jYJPCP/3GnKaNOpY3xvHhQC/5AfoCjhnhNG25jtNcNuOHCvPYv/uvmPf6/ikEZBJx9akUKg8RhyE
50QHsxJb5Qo2S+gUA/QtZxnqXy+NGU1kpEEv00M1A3YJu6X9RYWmu0oZbXZd5v+tevaUm0c1LGPU
OF6THPinO5ubZ5SmqS+dJltgtGNaetELfPxmOOW0Hg6GjZWr7/jM7mw+1L5vtYrOJebQfrFd3Lq8
oCIboJENUWgD/PNKW+/3kPo4zyDmIvy8P/TegQ55Jrs6ilrBjb1PnJFkK+/DR1/wvRBYznOIBcnE
6Jg4OHmxI8rqvD9acDtNuhgiuRn0Kv/sgR58OdTypr/8gsjfRxV1vmoYwK4aONU1UET/skI3jvc3
yhfe5PyiVAE3wsZ0nByVfHiWD6NL297XcrRgcWg/AE0p4hMaSk7kv8h8qZdxi/zuntIOnrSHJM23
PdVQgJYgjn5/YKeO/M/GbudlUibGxrjc921Gowode6TxgiXw4whuNcW0uayJUFjZjSiC3puEHstX
KkirfagDacWL4ZNZl0Aub+N1rrgl785Y+7qaWXDZDaKANcGVyrvDWJanjLiciaIDYvI4phpKNNT0
1fezPn+LnYb7dL2Oe8HIaR8yrdLB1NVIJEa9ISrOMwHVVH14yD5S5i1iuXk20AP/+NJ6hHcdwoES
Hnp9wnmL5S5Ctr2lKPGMwUWLke6KMO2E7gYKrWR3fpajB0KyTsjP/WDI/95mXV4U7pdOMonKCTGW
VxVT2rWh+81BLMfP6B2DA3x9GTk+tI01oT6LP/R/sn3VQMO5vfqVPDV0OAhLpuxJIWG8E323W8O/
sLyGlVq/r7E7hR01IccM6Juo0Irptp/U/KuYU0GSk67S236qk8p6fpUXJXMa8H9/b9zHN5z31jzs
WdUHeg0hmB8AIedoBjglVb87iAs026LCxwUzOdjIHZ6SFNUP7NNFgVdHGE6Mind0+sv3LVGAgMhN
BIZE01h0Nio9qOdnrJGpOtSjlKDpb6eAldxI+C5O5tSKPbKpFgp06GtisKe8Kx0Ucnp9uD9NjZt0
ro2XvqjcBM+PT+kY8ukevBkfFx9OUsaFi+pYXbXjaWY+1QU08wVMiSIkrAZ5JiOpXE9EjVsP3+T1
EZ6cvLKkqulMNjQq5jNpWO1ZSiEOQ6zPz3Fnm1Ne8FuNF1eEFkj2Ou7fq/voIqJYoAyBZRquMPsg
hXLagfg/U/tyn22UWxrRUY8wzWDcTaKQoBrINgUn+RZmpg4pfrdCkfBwDXsoWcz2GziHnt4nH6t/
sv2xdbec7laiGIW1W9KZIXGYSSDYkOKuOp0QIj0tzl1D+FJi8YmJC3mP5vbPfQsTSUqm4b4G+Onf
Dl+Fm92zzQ5VOMDEP6rpPvayy1wckLn/iLbktZkIjJvUR6BW4Wl5lxBAJST5vs/O0cty1mArbzt3
q8UlJYTOgGngD22qBSeLuH8qoYSpg/VziI+fMKrA/gfsHbK/QP0U4hQ2zz7+HjJkvv+8WNytaWDj
qtk2xgF2DoX2bGqc8DtrKcH7CmxqBfxliuLgHLfuDk1N2tNCAnGr3RqWJw/m+ijauItYwWrKHqaB
184aWy35iGvHn7ufqo1QMvYvov9Ak5B6lP0Ke1um+u5cRjfIMht3dxrIiniCfXO+gNTZ8UT9tDoN
onFMJeArFLdRPDLcrTRFoGLk/JwcMAzY+RMl84yEySZZ1Nn59JbL2/aLhuwaPeTn/+jmO1nhuJTB
fpfVpCY/8ZLSV14xZqhImK5PiK83lgnkissEyp5vQSIexv8UiZecvUM0AGkh5HKWoe0x0f0rdufW
+eyIvZCkVzBssdLgyTvDsY+mY++eRJG8p6Jeu4YHoMvBNq2pVBpacLJwEI9EqFoe90zR03/KNeGU
h7kfSLn2vCb9n9XAcQ+gDnjXM3MepFR2d15/IC+1bEvws4Ap/+vjaENAj/v0Oji8Fdx8++OLQYzE
CVYVB8tNe/h8wYflDBGKif4ZazaTH1oRY2GfPtziV3USlq8hK4F4VGps6Mf4hPqrp3JZqjcAoOX3
TpnbtwnqJr/7BNFGSG23KZfs7X57w7Bn8WnzoAxQ2nJDUtUwK6nHNUYsiFp/efp06OBJy7i+K5N4
a17SBi31aWt87YCWRYtv4dC2ZvoSkmzRW3b91Epk23LmxwKjGZXa7yP/C1sLaXOXMOPWY9tBiOU9
FhRli5QQRIY/Qg0QHyUaJp+Gdk+Gbj2n2Ah0wgTGkaaioiP3oy6aH6rA/0/oDYSes4ONlBDRnRhY
unSQvB9IfY74kkSNnuZackMD97nhXTahJd5k9G2sXXie0p7IZgogxQ+89lMe9t3Y39qcNJZFU+Co
VInStw56nMr1Ti1PaIFgLGpoUVCzYwTGtE/eeljBlwh/2qDKPf6WSp7IkcOOjS2KvSD1Yyaf7r5g
kisiM0VQRFYTXE32QYu9Q49MJUPRkwJ4gS5YU+StXttjcs/s89o/Cpy1nuC4qFeQ37WkRpyYXTKk
tLdYGhsfq1ZQDJ9R2xmHiQW0k9KCJgYoNsgdp9SzJIuv4BTV8FMBKMgiy7TkZ4XEQkaUYL7AQn3N
i3dAxvz/kaeG2q+QAPIkGcElrALrfAmEhzj4oLQ/FZ0luug6KRm1oZA8p9b4xrjgRHtDkkits1j0
N/IAmwnrnqDeC2ChIjJd5O5YtS0Xe2altiSmL2FjCuZGKEc3gA1s/i2uqt7QBbDKeF1jhUYkYKAc
uaVFatT3ik5OgypwzoyomU4zy5QGZFJLUbV0so7ykSqXdJi5ILehQZwbBX1jQKNh0Fi6t8pJDjw/
NZy+zDHyykQ0TQS+0cBoppfi+FuHzqC04+b10Fo0CrOT9KsEiVeHzVou5og1DKcSUM9QorN1Heck
FqqHDYay7FfeObikQ4nb+/4d7cSvQ9aV/zIh4OkM6IdbaVDcFWtXtxLkCQ92q+Hi149QOw6312+U
AXpDLVAtqilix1rXaMfE0IK0r9uwLBf6C+Dh+vQRt0jKEGztciNuaFA4/ITCip0q/ElZz/ivplym
w6dVlTXVE6QmUV7vnWnqFcOFs977y/7Xwt6z1bNE8ZLl5ua4CHw1fyMqzmABteO+fW7UOjcRAbEe
z9BCUGk85UEZiQNJG3uFMGzjgT/MgmY9WElDY6eEAxZthp7xEsi11r78T6Lxla0kBMeITiTZxHcx
1bCdm4hQcv2gcMbUk/AuXqKs3tBmDOaG40CwtAwi3OddihWeHgkSIQICcbq5oAZhJbIUVZRhMUNe
9NRK73cWpn96peNolknhxaCgjidAopJvzhdSYRe5cnIkiUMeut+Tcq6ovaqrbQqM2dokDwY8QiU5
Uv6KyO/c7ZnICM117siGzr1ML6np+7ynSn1NLc0T3+gdMXPa/SUTLJeZhd1QOHZmK6Z+5XI4LViU
pusTUMiBX+14YEYFHdaZkX4PsHK4oaTD8Z2y+mTe5qM/a2XX8V3YE6Pz7Cpbdj2HzcLNKwAj5Btn
HVUe5zVlQZNjmGChycDYVmv+0m8cuH+s70PPkLreB3FutLZkHbVmwvyXqkLo9mAYBb6KWoKyAQ+p
mM9Pewb3VqbjLsgaElBRPo5+1jzpMBHQoL7x18SOWD/wi2BLfKGJJvAHhlppSpvx8BdZheXGyy0/
breA4venP2zdmC9SLK/I/lcJRcwy3ypYSCSiRlfG/fH6AvnBtd7hXV4GuCO4lgEOlh98xiwBhkTD
cf1K41MWisVuN8zWnWtr/L/zTNrjFjVhgjeozNqpWNAsAVAXHbkym0z3XCT6SG51OiteCOicEGmb
yay9+mstHezFlAwv9hmuwBXTHUfP5VuKABd7HIsyk8NW4DSfGkUqoRRxH1Y6loBS7QuH1z7IJrsc
9kvRUMQLYtBvbzHDH+SmrQxYrDZp8g1Qb7pm5P4YWUats7v90fNWoiIfvQEgqDQaP/ATMIecUCck
mZ40sfGiXaH4a/ymDyKdDSDE3E1J7x3+OIBhfxHMFSCsUT4g1dtwFK2tvyDKyPwR3SkxbucKRuYo
Lx8qb1aPYdKj1ALKbzbrx3OrCpc9yWYkbp21xJ5Ue/rcQfPu5k5o1tyIAJibMCe+gHVMfsqwktpp
5rDfKaQB2pmX/8Ep5zC4+nrgwJf9UYRmDqWfMOUlasJ6s8yfiZ057gKPi1Svwft6+6pOuRLA4kwz
WPC/7PvkyTktijmx2eAmYw7dUtvK3MQ3z+v+jyWSrX67Zwq1goRCJCWmEY1ZTeYnZ3kgJGzb/Sdr
HtrSNxHA9WRydY1z1KrgvmgIodRzYnpoaCOHIoPWr0IM+z+MwDvJ5uErxqFIhsOwL4xU7/TDP/p4
9lvQm6AG4m+Gh6VsDh+M4+2lKTzi1e1m75RA2jtiCalI5bdHVetFJt+XX/9JBmcktZqsgEjHKip6
BaZhWNSHebJwtmVqGDiSb5Kpc2dbfi08cp+dZKNqZFTn7gSwe0Ir8laLodwbtEyzQSWJC5sfieVG
eELsLgy+L7vWnVpZbAqov0Ho1Z7ax9cPokc1Wuk+0CTeTedSDAkj6dlI/KGrd3D1uCzIyo7Cq2NA
9Xq4Tikpyw2w7OO8DDJpSzbGSpix4uW6SvHr2fzhHl7xdFruJ2mnM4iOd15gixfbVraNUFdfs/BP
Sgfbv8c0TCizzm/0c7cQdoGut/AqFJHWZqnfxLKvZyvpIOjvRkG4BAUTvES7RXrMz26wUVfjw8p4
U4FWQd2PSLTfRcR3JKwhI9QGpQbI7niBN+exXgBOdjp1YaXGVx5UNWEXh7Qx6SWGbUHPtChVrJHk
HpgQH43PbxSN3w5pPYvAEnOwBrJ+dDyEbeOuzx4ofXG5jrUevPoNch46DLm86CsfWwcm/VqZzKOX
2FZLm/FX9CVUf/eGg6HtYf5Tj7Gd9AGAJc3XNa9Nv9qD2dFKjsaZO2ZrZ7dU83spmj2Ip/DpEdq0
iZQR+7CYdgXl44KjReqJEOhMsW4+4bEITpRMKbHTOmpqyIwLtkNNiiJOA0N05KyAtqd5Qj+tX/pv
zA9Uoub28yJNoGuQd8bb6l7XBXin17WDMwL6dlrlG2Q5g2m1fkYpgy9Gp6sGgwD0z5FsQu47YpC2
2W1QLid27+pi737uv1V0k3aMWpwTwQE/7TGsF43migYZme24CSHcbWvPnAniuJNPqr8ltuvDFEJ+
mdiRdrUahEQG6raZ3dLxP2NMJ0D8VKMn9FfnHKHEllwBrOHiEmR08ZgvLmHVF7FzGp/hwb9lQxql
i6CjRv5rNLHQziGgg/gfUkbvDr/KA3sOYufK9/s0bIIgfOfQiugVdu46vKry4ZBvGCs23z6Tr6z9
+ftV5tHn8qZRp4uVAaLy/9dY3TClc1EOYBZWbW4wUph0TZpvf7VTUEZFs+U3xdrgNYhsh9PZUFNX
I4YjIwLyUJNOWIBR53h6WfwQkCz3ZfVUYzxkkW2r7csA7r0zH3hC9l9Vk+1CWK7D40UUdYl+DRsB
x2QkyNC2rDdqyVdGsoupmTMHOkCRkZOpivJ2fT0SpE4WEPpyHVywDXu45BylJPf8NWuSCmaBYcE9
jrrlViVN54geEAP1jmW5355FjoKTGq5sXnHWHfY6i+xPeJhei/b2ofRijxFhIA7FuBpGqfz3+sl/
pzwmMY2N5YXcTVlMep/PhzE5DeZrxRfogXnYdvkOktyx1wWM9aWi1SrqB3e6mZ95L7/7QoHd7CYX
l+qq6pQpOubYJCQnTfRKIlXypGgm7nZvUGKpH6av4yZJ0AmkM38bBVBbdqC5R7hPhYnxEsUAu8fi
9varg/BJ6zj+PuYTv0/OghitLtv3i5yUHxgfcdIKeFeuBquGIkO99qA8+V9Y0K5H25SfAIaswnq2
OJ+99sYo5IeopElCJBdgwtT/Em19bWs4u/nMwcWCHHQBolnzeACbY0r8oKyHi1T97UxwTdGtweO0
vlk+oKAhwEi/d4izod3Wh0hfymV44VGWaE/0gWBT1pLvyYum6T3PuguNyZ7ws0lsstBvdZVF2WQm
FKKQa8b/FVW8ty2ep27lCdDCY7zDrak2aZXXNJwYHl+D9AzWAvds03WqQbM23oLG+kAne09RT3Ro
Vs3oaynXaJjSANpfblP8NEAw146KlRmPIWKxE5yfFMdfdUp+kNz9lVzYNJSwFNGtLyaukvuEhU0k
4XYy8N9Ei6IdNBMPN9bK/U6O6y6Ze5QhN6ISsf5hriUc5LswEdZIXgAh4zkC1U9J71Z7UUom+d13
dtTi2Bo2wOsi2g+VsZpg9SZNH098+7zXQTBvgk0xl5I6u/MzMBQwaCm2ix6Jo2M2Nf+QVMy6bqnT
T8UdMUe9dHTmi/pA/EXqKX2kJ+HKnfV5qN4VXkSXiylFyf2tc7eSrS/QH6mML0trLIdR3ssxuw5x
bErfwTW2qFr9W74UhHlhEAvg/x6foktCWX7HNO2M5sK+yq3a431H6BXTdj4rOJK01Ov/tt6R0cNu
ZmCOsBnicyy9v2LhNpfa2EmInU/2Qej3ZSvcON84BG/OqrXym+D3NCRaWGa99zsZjChQKMmhaHxB
2w/Z1UN8qZJoa0EMgquecgj9+6hM9plWt6kjIAMz4sSuMw/e5ihq46hq72W5UFoyEBToD767FiO2
frHc4KtsJlE08a67wtTWVaW+gZkoQmSLGLODkd5fXyib0wiI8DtbnOTu2xxubmKVdf4shk6+GACD
nC4lyzGxGaWQkubLKv9TQsFd31R7V7bkgAg3wexm071cNKNu3aDfht5EAoJwJyCL438/feVVLJGu
yIrLGkGPM1pl+7at6S3Ak57dyrNDGt9s3FlLdtnpc4yZwYJRDlF3odPB1lifDeM/ENRDqlVgJdKP
zoKQknhwo4G7lP875s8T72rwoZ2dNqdCgD8Q/yOY8kQeVNHAdE+OYYJzOLz7bVMB5n9Saz4DJ/4n
dK3o1Q4UPP+IL4slKjKRd4nQHgokjb/tS0/Y6RJLt41bsyGDwWe9Ws0DvsXwXsahjybNF7rh2aVG
PIu2Jcy7LaMnPC0VzkJ5SyU9VJ5737CD9LIiGlIFZibeV1nYyBWXTN8AsMXuhtUGj8CPaguGBRn3
cxlL03JPniu9ETGHy8IfXx6JdXq3JWExwKvbk/znbO+Ty/g1eDF/4Y9jBHug/RIoet8YoGJ1r0h2
cm2WZPfngkBjIOdcZVhJF0wiCceucZisAyCHPCYGffNC8Noaqk07iYzUDTOb4vMHJ2d71Z3rQCQK
4WAuOlPAmeevhDhb3j7zY0H4bF41PcaVeOJgZgULxucL2R4nRkKp/oezvtqP3AOK804N9Y+pJEFZ
x95HpPDdbrNiAETOtMvog0PMdbyJEl33VW4NZtUxHz7xYUn1poSYqB9fJGr0H8zIy/KC8b1sqvyk
ai5WM2ifha/egNwYDOJOIWloDHR10HIUeREalEbJ7UB7ORt4Gakvd4LAwP53I+xdWMZZcYamVI5P
KdcO4/8RdkJnusWRrG+HMouc141wHjHf2aNmYpNOZo/yVWT0zk56ZXpQW72y/QIs/zbHrmxSgtJB
u5JfMQTXIKyWYpNB8DuLO81OdyXiUbjnrHGqg2oCXEBgfj9aiGPTqQ7Zf0NxpY9s7ShVqqcMCOpB
5SYTZVV97baYXSi6eVfCAfSUpfsTPlWrzTQQeZsdTlBIDuOMS1TWXcX9PBKB1gra7EWGwgWGNJwZ
Tr1tYur1ndZ/mLJewZ94W8Z1y1xmSgxtGNby9G/6WNLubBF1uBzR/YZ2z/dP71aTUq+OKf/smH5V
/0UrZe2A03lTNjtcbGXV4Dc0IIO81ITqIb3J2kzyRx6WBNiEULwGUFFw4gi9GArhhjqH1ZZjn6mh
Un99BFQNJ5PFRXlTkwalGO6ZR1GIfjdiS7PkIbxCo+d41DDkQ90Kwkb6wyoNmfFX2LdWYfqeCRxj
yTlYin96WndLjioC8dsQV1cghzM2FA8jXZz7M/twpUrCoygJCXYdaYR1koWyl1nH8oQfz5tDrj2V
ek8NPR0AvMTt0pXAUiqfmYdtI5CPiNBQO1LEsU9hgrQ7IUDgELuxkTJLXLN/PN8PYmA4KTCQPav5
9EgA3CTqEd5atkeSOopeYC/XLK4/K75tJXrhU8wMwq01DkSpfK19N6hMULqVnJi8TQRTqanvWfiQ
IrwjSx/JT20hN/8tw/cehDKAQlQaYsZ50hjXuKNReE68kFtXZxKJ5hesPFLDjJhn0usFawpniMDk
29mxMj68NI48g68Zs9wyNKaybX7/UmncmTA9bFt8QXGz1P4Xb+rZTt5xP/K0XVdPO/oJEN3R/65d
X4ZIQybPL5kDjg12V3RqliD4rTfRW4fhLHoFH1WGfXqqQfUJS3umHkjs1LLN6RPVXw+4AvT/HJHN
T4zfR73v+VV7DZZyajMZ7p/a2HcTB7NpyTlkLKRbMxkjHz0US4soDVfO/z4XthIwhFhKulImdhL5
wAaTPrLhdkll0OSwg+S/TLMIz2835jGmN2sWz1jbmGQwy841Em+jP/te/nKZMScUV18yEwJTjGSs
CMngK+XFDPeIXfP83z5J/3tNv6V+4RGBQXgaq0HPWoq2ARKzmE6lqb4tb16cc0GO+1Aqj75ZkaXp
zG6DP4DBGSdhKBDlbFGnuREt1rGvFeY98BUJlpacwQZlyIy0SSGyLHyb0AA4MhcZiqK6UH0YT/wF
gGF9TR7dnzjkDSJI/nsZaxOSbJsc98bVQEk1bG8kKB4FwTtxozKlk+7Y+fE0grvhpw2dSslTySXQ
ri0gP1rdZ2xGcIdSDJ7ckI8XkmsyRP1evlQUedmfMsoQWOq5YqNRD4IguTrZipdFQ7SEMonI79+b
pIXpXV6eL/yNZgKMyNLnaneRo1M8CdY11Kh4lyZc5uCaT4Ho5d3XUHoahQ+8IKtmxSEnARTiV3et
iss8sKazhWfh3SA0anYCoEz2Qi7MSNjMuaDC7mEpnoaI/KFpsNBiJL1DG5i3wqoamLigcQRtXvvh
2NNMZ5ZbADCaBdgig1tUMm/rVE+RZ6CZui/XnpxrSrjq1NNGJIjEEPEdnbJb2GR0MO/KzT3VgNwp
TYk9bJK2qMrXm+AWExS6OPqgwKNBy69O0I6/uCANP8yZWp0IL2R7F3g0/HwJmq4EQGFLo+zr4ZRw
RlgGc3fIk/iApMBPsBVaj8hceO2kaCDJi5aWzZt+1sA3GBHyc0D2HtZiLwvpkaDf6vnEL3uSUgyl
X32BFWrROIh4tbN3mCk0XW9+nEyA6RxXKTMSVcdOlcBKeOkZJfH3c+yml6BwEDOfB9hbvj7So8uL
qdDiL/Nr6Aj/1bWhDqHWZB8hkcZgthDTZ+hbazNcuB1bjJ/MOcbuffXdWuMsf8aqLN9vvs+b3BMF
Sobs7x5k8Z/piWih3knkwDiOwjvpF6womz2nAtwFqakjf819O2bHvEe9/YdJAUs4BE3X+PviQI9v
/bg2IyWc20TY86MIkTizihdgRonjqYKKP1hYUjkr+91O0mvv2Bbr0pCPwQzOyCJOp+ayuB3097h5
ZeqH2mL2axau3YHCy2MOoDqXu+HPWwoLfSD1dthCkPsevlE1vIrrPOIbBlhPq5WsEb/g+RdRHq+V
AUS/jpnvAGP4cnJVr7VaYt3/l0yBgfyVOLYYIka3KS7QxVQZnQDPbOEqucQ11vmU9+anvdslZHqP
tJe/TjLI0N1RmSpFt6hL96F96IfeDLD52mWZMWmaoouN5eo+IYBYKjzcjY936JoeaubpC9U4jai7
Hhz0Q/bDW4PJqOGC/4cF2lS77LqX59qH7pznZizlArmrq+X6EteKT9NtHrnjqBqY3FTvnmNGz441
/IlNk9nFa4VAR8rES/mBRcLR0zsbp/TqiOmu8tPKk97TexYUQZyejvZeP2CDoQ/RVb1ZDOuIaSYs
V4K/LWwmLwx+ezirR4+5MpB1Aupg6zZCL/ehvCkLIU7+kENxo8ndfopdJrh02qySZEy9KHh6sjET
A+RoLQBnrIupOg4G4uP6IS7Ex7BpYaupWGZPvsoJNWkegiRog0Q6FS7f5qJ2YUZ8zbbsYpwIDv9b
hxZ8wjk70xD0v2zioXAdBl1kHRCU+jFaw4ASRJdxiPMnFZ8+TT+NlxBFRfqpi1LKywY7bYj4ePZK
z1LM5CP/vNydehwa3UQzifpB3VLRxfSVrp68LOmcmXe3L2bkjeVRsKWiYBJESUsSsHQIlPbTTE71
BevhWdEjRoVmmbRcNZTaZdgHnBlcH88xR+1kbmo/n4Ig5bMHEwZYKqZQUOt+Wg73T6sJOi4HKSkI
J+/AYJblU1+WjEJOCwWo2jTWpdD3jNGTwE3d43zJYFWRlON3i6KOXI8miSDTfchvWycNLngAV5MT
WBXxov5Yv65u4L5XMqgFNFfIwniptmLK+mPPe5+/9hVK5JF2wI5rqSx6bYPMkeH1iEjTkAgsg5Ao
MWD/qwD49OGClk0Bq7NbwvxarkUytEtJbSLQCR9w19Kqf9CbL2+VOb2WMRjhDW22cNrgpLiWtJrr
PNheoSUaqS3o9/O9HuMyXDrA1MwP+exYZq00YodEFGFVdrkhCNgcYrfbh5VhjIXmRoVfNTFkUKDp
CfwjKykdED4aYrHYDA9r7rAcG7rZW42LCyNlEy6Ojgk3/hfmUwGn8xjuM/BD76tbthfd/IyX09Lf
Z8vCp/2vCDRykLN4ASspuq5e4PNM3wkYCPym+f8vN+m/BfJkb9q5NqDOwrTTzmbyPcDsbdk6urWv
qPGvBrGHhO6pIUDXvoYjcLt3/HAFgPMIxJkxnCCCmmjyfNBWYsPc0a+e6SRGRlq/iF7GiY8MR4zX
gQ8Xl1bRvsSV/ZLNy3UwB66TpnIEt90j1XTW+h0HeufQWoqgGt7TW/5j4XDEDaEmhVAlh0x69a9j
0Kx3nYmIQu08XIjjeg2TfsBzyQMKEkjzjBH9d/Sr05XGCplMfFt7Gkab7j454IPi9MvAjUsTJegx
agmDdbpwRm7VBu+M8R1zqEJ2wNRK0DqhQ8E4xA8AjX2DaWanr5s9l0a3LRmXuwiykvOa8HpAgm7r
z8R+WI1V89BMS+afBvaxGjqIfjy3/pUDqiPq0R9Z1M2k64EulmWKQth6GdG6GnbnwsC+tGq6z5Il
A8lVL+QdxWk4rfQeYjEJbJB9FUiY9thdv/GMkazhLGunSYSi93qj6yY4TrvSrmvDtZEr08dXCfM2
HjVAZImTBZ9I/7b045W4pfJ7EvkqSaLV8LQJY6vZQ6SywtLIEc00yOQdxMhxsEd7JYbN4eZTJGhF
91BR2+8sGXjaXOyzcKf2WQMk0nqHl7jhZqqBKEdhcqPDIXY1D8Vv8dQNvLprxTKcUZ6FAf9mWSS8
DNtK2swSFBUjkYGFWBWR0a+JyJqFg086odyakFmgt3NC6iQ+xMj9XCjhwxk7DnufiVeRdhSqRE2r
XMfjKc1u/2KVDAwtbgkhDPQMsKiTeJKjvM+ZkvnShixfjQJ4qgCMnBACXUC2Hi/CYUO4Q5Mcvsjd
yBp0Zdx66p5StfF7FXbB8EBDUhFqAqNbn20jC09WFeYrf9XarySQASLXkGp1dJH1ZLVleOmuEkdX
mzWcjQYx/tjQ5pm/iIdmsvfrFZWZs7fXoDkvB+5vkcS6TwWoxdbhmeFQIj8i5n2R04qIgXEE1Psg
8TW54YZJ962f1jY/t+Pb/vqNiMY3ch/MNktbEP5Na9TrBqh08CF2JZDu/7X+Qo0Qt975PUvc1XI3
4sO8rn2P31C9sE/7hqUYtBCb3TDtEfvZcOAptcBp2wKW2P0oQIOPG70srjIyER56Y7q0ogCRDD/x
O4bjVVAyXip6wQIUJ1nT7mvtybG3w+o/zTFkz2rLGZm5cdtDBf1ULrokdW9FIcUGTNwkmYHT+U6S
cCTNoMEGa6882wiGJMx9RrmlyH3nQmwuMTMkCgMd+fsWs3eQvUVAGtyLii+Fs3pxx9H1+Ve/Wj1Y
ziPJtDgY/hLR05PdTuWvKdscUtTl0ekt8yiNakjUfnWes6Sg73+4foViTwP9jZ/JEMwtncI1UZ4n
YjmRCgBO2tbut/lBxUTeGcVzOD5Fs9KSw+6DIS/l4iPKA/mB9Lzt2FtEqjReeonjizWaJkkiopEN
ev2+JTpTlnhhDXaExN8ZBLQBX1gp6n5bGHTBQQF3TmGGnmYa9T6FnWyzk1iZfDqm2AyBLt0B6scU
YrQi5mXUioXTeiFm0D1Y2zQcnG5VbtL+Pgxf9jT7iyKl70Bp+gVYDNC8Y4G0IMLbWdbWqyNiQTNn
JJSk/0hn4gmvqDknim+LkYq7R0Mxl7s8Nk5fK9BVjsbDlXSh2YENXagCfC6QBVM+yBlwMyVukHqj
j/E+ujZrXZ8jY3rqgtKGhbTfjSaWLJtD0okfQSK0vTfG3+vvndJKNyjl7lpOPKR1uiaUyBrYAYdu
HZAkYzsajkDkbKQ0Yod++12/zfPI5AUxxp05FB/+ta3rEVpOPp9+D/m+FSyLSS3KvMyuH47CrXR+
3e7jDRPDImicg4LskO/HHJlK863iuEuN45wuQx5JmNb+SeXQOtu7PqH/0fiH05EN87KSTrbBR0tN
AkJRWDzaaZkym4674fDuSCqeVnp2D+Z/CG9UnE7+SItcLZSiMd0wbFybrpO4qMVDPNcbfOG+XIR6
8X/VCh7j4hGuksBdsRr/jPyQR50PRfZ/1giBSu7J7O4LM5bQGDqQd/Hvluh7934uUjQ1YqFnZMWp
WDO+lMlz6FH1lNGuX64tCbQJS2eWGhcwGTLZ50zOgziW+lkrwiKKB3rOEfaAcwGrVPEwmcBVkZR2
m7spp5G2gdfitKwh/yTmypRVlgfc+vCynLuHoszWHBkk0IZiAzDkz6PNwM70HTTqSN1ztKAy3JwE
T8p/aSfGBkJ795X5z7/uBVV3JC4S+qSVIS6NGq9zIrHPUs7g72VADEjna/EF+vOFmzl73OlHy7TJ
jRzRCj+rw4Qwnp8H3J4DsHekNZ9i0+l/j2gP++h57RoC+LG0/UsvrsyXKyg0XvT2vm2MP+LKEzb7
3Zh8qUuq9tf2oXnIAQJ0Ak0f/LNpeokT51Irn993r6Z2Jco6/HQOfOMBhNRCPu3DCqW8Wb1IuD5s
0Xu4053VQNnw0AlQR/Rsu3rcKhcqzVnNKQUt7/EYa9qfhJ+AbQPC23tJ5wRLON76KCiNure7zF6S
AAHw+Olc+2rEcNZkjTgBwLkm/9DbcZj2Qu2HJvQNesF6Uh5rtT0oU2yoxqfhLbGzFsln3o8PrcYw
hctSQWI/NgeC/6mQQiz3K8MdhVyTHKaBYrUrudLhJCv5B99t0PnNCqUak6qtBKygtXMbp5bs7fcd
hT/2qI6jUnxAmlpBD9GXM4zZf6LBttktiPOm1hRS0UdsvQ7N7wVDegv+BsjJShQ5lKdgH5FkD5FC
gnLr78ouFa2a81Rrd4UjvNGYJLCaIFu797CrfE8zDpIXCfPvNFJ/3MPNgFNAEglO2CmXZ4TvkAEr
BgVkX4kyCG7Z4SECtx156gz5PZ8Fq0paDUfWHOSze7MYfJzBZU1N3OUGsxvG2zF7zdMu0hQjsxG0
OTXgqEbTr+Mf9dISSSFxirChlKMwBNIL7xWk5fR5eFJUT8xAGIZKHLxgqmVw2aYr35A19pM8HBGM
1WgJXKS3rrDicFVTL8oA0kgqJKAtK1OdtAMTgMrb7P3fu67LwfxdS/1b5Wb24aLr45CEzPnq38vD
94YC3QMBZGkxYH5ZWoZH3jIll/Ol45fjnDgRNG0h9JezYlYreR7bmv6Fs/8RVWVMj3EWPS19m/E2
urGm
`protect end_protected
