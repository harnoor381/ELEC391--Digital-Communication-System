-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
ZAGFrZyY9cEpzuSLUrIKehtnhImXaRIA/5/Kyz80awlq2uVIFBYuDiv9W5cULnVI9O8G1qc8GBdT
yGndekQ0sEI3cghHz5ji1nq+5UTENgVJMyKOrKuRTl8wcAD8jzwoOOiEEB1LwyDTx+XNT5a7mxoW
vBuN2x/gGKY02X+nFczWrYO6URk+V1S4BvUo3gIrmbDlQThNUqd9kLjVhJauJua1JEbvWNKj/bk3
TxmxJjVJegBeVobw9r7108qseknHTou2jBxBrDHu65rkdsJkXRSmhQQpiJ++2hUcDV6MQBr+COM/
Cldjlisl8eBtfg7kBlfo/MfA1GWdc5dYio3kXQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 30464)
`protect data_block
Ti+vYyRFpOiJGORqNeCQdoTX/8qPNkXK4ck+plkZKVMYYb/o6/3T/+H4POy2YrUhR8TXVKSSrR41
XWubatB6SGavkeeHmhuPjI6JSOOy03vLRE969swz3fwpB0P//T/FuC0LGKuPrtRLZGuGgxxDwyK8
uODsDOqGGJXiVX7oCDTQTN/CaiZI9pBeHHszSp1jSY9NRFqK2xwt6nrHUhp+TdBDww32aX2kW96T
Dxyw3QYmsLUMc5pDTtKBkwHMzgCvRS2ItQ5kkTMNKE6ZcMuaLovRHhksM8tGZE/p0lOJQpgJC7Xt
6fJvMONxQX5iGXHAH/1YxjmxMAQCHZtCpVdcPr4+tiXzs99KMX3lwPnZwI2m28+lyCu8lRPYbwyF
gXmDxJb/dmoNv72brPmeqTPLP87ZZCmxUFGQ02txkcrVf6Tjhe+2GRZcJAFzK7YIS36T/P9Bs/8w
ybngx8AuBNY5WBvJxvtO9URZlqXZEZjS82Dp23dDAyvDn4aGTB9U3+VC6Txk0wYT7vg5EaK6fx2R
sXuIkxoYDtl1JSODlqSXdjI1YnKpNOT1Aqa+Q3aavPgS01ccr95WhyG+rmkqm0o+Qf/EFSXqSyd7
KVShkTWRHrmUPoDtIL0CusLPk3wldzS/cVQsuYsXoL1VvDosrdyaa+ekEISQ47CJu/UvGozxOHp6
xQAuK91FphMUq7JkuTZGklad+KxNmrEivEIBCYkF3HUDwBWlU/JKV/tCfUnpC1Bt78NJv2RRXQMG
yiRtbqhKHrDFa1yQfiC6Q0ZFBLJ0hHstA5NXKSWXl1+MKP70nbcE6akgpUWJghuBlwsDgPoKYOIe
8R505rujsq6fJE9Eawl10sfEsP35KzzpMI/3Fft1U5NvRjczBfFPkaLz2f4AVY+BjqN00BuRsUmn
1u/JdOuHy/SUXf05U1uBT1UFYKZOPGq7Xtlf8HKk3wztByXepv8+gKAlCDWDdzxohc1BFp697TqO
47sm/F1XnmjMBwhM1MZvjPaCSvJqOBoPID+WHzdZ/RXYABJm/A1wVr7RFH0sl12xJkju1pS/EIjP
SrG6845N3MLYtx8IIJ/Kx5qQiSLalc2x6zD2B8yuUQhIzopjvEYCbEjYnjN46ol5K6rdijBpwEC8
Yn/03iFIQ4mxrlM1TuBMGNmEjChHSmsJO07/Bdb8quJQ/I/HzeXZ1eLMHsWxcOfVuxywCeS18jNo
3TkUDAqqH296OIdj1VIp7N04H2mrQZNFLBI1dPfdJfFWJ/iprZm0xT+meN46pyqe8EXij6V2OOn/
AkITLHlWXDI5MA7GVOPG74FwZlblbqaz5AMu/BIyWlGFCjx13i31G390RQXJPS1a/TDjutaI8mgY
LtETUiIY2rP67TXmxy+aCem72msaflNsCcJRF0U8Nz+tWjkjw8hUjI2Ld1YFn8E7r20xHW+gZ0UL
gmxVrbJxbpuuem49+8L/Zxcn/hjvpsvoRn+sxIhiy0p1CXEvKkArBYR9t+VNm6iMtDy8I+rTp6yj
g49/hVrFSaMB2lCEf4J48vr+nZk9hhPKXm/xzoQP8plVzeKq61lzIVKJd8J3Q4O9Hiq7F/NoJeez
vVv1ypGZ6XcrCyEGnj88bHrCB2Ja6as7iFoAot0QMRaJtwwi6+LXhUjW98siYXywJXXDbV82qg+P
yQlpLaXPWbQpZaVZBHIFcf+LktqSsLD6MzivEhFRnDOJ9RgKsFGGRwAZUmTJBfICsejcLy+bcABq
C3f53qrjElvS+5vvhPlKgV5+P1rFTX0M8j5ZwALKrk6UZKdnzO5JVpXNY5OUjaDPngB42SHGlbi2
5kHTQX0vAtFcLphOyZtbDvtDEcgGgTaRkHoNHv7UwXsvgpW/OG4FZcK3XeQiENUdVeCfxOve6Hzi
w6iZZ04hagXkQdWi99IS3P59n6qOQY0vq6p11Mmyi08a1nzWhVe4CnHAcwW5+QMZx5ULGdxT3Nml
L9V6i7e1xsgFFsTmJ3dCHRlaELy5aE5tUzOQ5CU0GBB3wwkIWIwJRBH1hVMl6t7hw89EdQys4W6E
HHMMaWDO2ycup3PuXCy52VLThA31jE8MINprWgR46dJimkxgY7I3Tzx/CJ+KvdMmdLjwB2ZUy3rt
uzdCR6LI5lOSPJLAAb1jHfz68qsB8zrsw3Qu8Nuy4TefXauuFgikmRigVv/LDheiPPQkmpCICSdh
svesZHmGsNe/vqmCa2f55kfo1PVCYq96lKJeuD8qHqiNd8+jevzJ0P8hdUc6KsdFCHg5eLVqw3sp
aQ+9BXbvTpC82HrTAPjPvvt5XRfcSqDpoTQLsZVLwdoCiGulZSkWAMOAJLp7NN3Da9tHIK/GjNlc
ksNCbXF5eBV5B5XOGwLLL781y3M7PHPF3/t4SOYyfQKiO/qUKC/NQO5Los5oTRe0MqMudzr1dKFM
y6MKy4ph8ZtGH0QPkkJhnqyDLz1gh15prKvNdkjprbyZJ24D2w/t15FFx7ZUtqRTGgqqRVY5kGYR
7qjJ5L9ti3gknnMOQatzRQfCpCgSm6wPJL7CLpFAmcGZ5N/vU1W3VGsvmyXnUjFvDu5TameaymMb
QIQVkTNg6VvheocdWQIe9OWGcbJka29M45FPMZeWdxJUmS07mOz7K/ck4qDDWbZwD4owyEFXAMW0
HnlfpmCCGgwKYqiyORQnkfdsqaV2qoRgd6T6QsCgYIzSYLjXY27T+xvsbun2QnKFOWJMvijuKffH
zvBi1LK6/N6zCv8k2/abSv1Y+hi2fCXgo7l/eHZpznvjN7r/P0cwhcgs3BiqgWjOKrLusSCF5c9A
HX1oI0/h7my+P1GPmbhfC9hAgddbU/7Ji0hY0dEV3IsNoC6u/pVzLfTYTaqnfimY25syqBddmMz1
c7yFkzZYLa6rlyIzw05QEA5ULQW1UItatXoOOafvQn/t8Oars9SlsP9e/HaBNZCM2x7wb7rX/NxG
bsmHTVU4MgaLgmRutXIwAtNDb1VmQwL/ym+H36UNzip3dcsjdJlZQt3EBK+EoH1j5h+zAkrjgJsn
lu7CUL8/i4gN14uVk6x3dO7j7VtY2sNYLD7uJtA6Z7G3PZm2uT5JhwBE6CoOavZmNMT+Gln5RNhe
35yHSvSmlElArzHxVpB0/t1CZjY1vJB3/kIqFLQ+wTGHGTHxTVl/rKXM8XQODjgz8RswvoT7PIcy
uJL3BcuTKnzSNBE5QcJ48f5RkOzQOqCdJzJzWCgTML29i9vHsZosaT/55RNJzGWzrrtf31e3ptET
W+lleXPL1V41dMqWO/e1BAbskSFjdlUIcJ3BkV2DUhGFm/h0TxrbREc4oZwwh/TMjYTkGgvE7Ni7
nq0/BPh7nZZRkloN+5nYsuxAKfrIL4spij7Ss2A4bd0dYuNwJCFyDklEUWzxkg4RtZxFUjeuVnrP
fuz32+6A6qzAmwdkGueZR6wirhonSTLnJ9ma4v105lcXO9umcKD71d0246/Yrt3n0DANC018YycL
RLPq5GAW7A0w0ieZqCC3RQ7ncZ67QqjlIeLMAtlDPfcXPvgrjRVfZCdjbNZ9TRLrUALDsZTw6G92
IcGeuh6v3EDLbBvW7gucFLIverDpnQjF3fRVm8gFYHWfNW6NbAoo3TSOCu/JMWt6zc5gwpIN6Erx
v1EJTik6zVpNigQWPk2+uZQL8OAF37KKfTbgcBu9b4E+HfGgMgZLxpmKz9bpaYa3gB90IsGRIuBX
PLjaWy7ozPOleUsWDiHOO7v+MZ76USPU8Ezjue3AJeuxvEbt3bbBeHWbehn/xB01tYLdLeZYo+rp
MvpH7HAauWwqDACUgjYG0X+GJBxNFqaEBDQJMiqdHHay9OKv0++2YQO84MzwrTz3JlaUYQogPx/3
85XdYzJa+jOB4ZhiQkoNGtKfm3BsvVK/OyW0xhxaNyfiWPPlGBiJjF4RStqkHbIQrzXT7IFZM54Z
2bAcdvODLIwouUhiyjL4Ct8Tm06dsf/n/D+HbJHlMeGYUJhJi5ydaJjF+cqkFtW0Vp5+JZTvqHGX
No/i8UH0m8B2Zc9v1+siTDEyuz6HdY1YIri43x1N9Q3KFr10G0JISZwD93nQ/41zHyer0lUg05Uc
gqpmJdRe3QygDpJYdAaC8GVI+lFrHZl+8oP1XwTYhPue0LGwIacoF3alExgNOLbnwx5BlZ/3xO+I
C4zCsorH+rN5JSjJ7L6Y4BXt8v9/tKM1CDaxFZkmUUKipwJsujDP9kd6Rg9oTHI9ItEm1Sv9jYgm
tv6FnOeUAYjwnbMdbP1WYBcvQvwQur/VCPeft684pmKnI9pSkP2jTvz0UXt73tPwDzArMt75XIFm
GBCdb9Okk0VW7F/oQ56NNMexiWZESgCkskQFm9YHHj5fAvmf7Za81plfop7l8nJTRcr+LoBqNAhY
Su/2EonfoJa/+/mLZnNOPVRVuf19Rpj5HHG+t0eqE7p9D7tqyHmYQHzUZXB+O33lUXzDzdkJBNT8
zRQO80uneEu9yj68sl9TRGJwTHxVzc21KOx7I370BpShAm9u6FSFuZB3wQ3/go49/WmHT8FC+Zmu
NLEp8VDdwhLgTipexGT3mBH5ONjlQN9kiCgmqGDLrL77al8a+2VGfLtMm7sxNviwrX4PpDydYh1D
jjN4JUTI36C2wiz55B7tYYbbZCmCR5/MMP9IVnISaTifzUDRe69HuUvHRn3WO+mgm2Mi8W0VLLWs
Qm1Qjmzlh+hv3FkEI3YVX7zyZ29CRJZ/Lr3jAT1rMNFQVY/U9KsyR3iGlvbdrKGeTp8tYec98utO
5+2YjV9Mr6AYwF+PwQZefoKpd3S/pwgJDNAIETwfdH1AUYPePsvPsbnlYCkkJTSHOQ+eYIcKvXqY
VBEjSlXTU0qkJ40vPCe86YGwlNZH3CCMhmUK/MEk/JemNCi0ho7/e0D0JZ1UkWJHZ2selV8Tv665
eXQNnF9ZbMQZFethCmnlOXGMYre+IuG1umll7J9Yk+wRnJ/W/P0QIhrS3W9J9xM+d+T55zA26+fY
bUfey4CsedRVtcAat3LsRvf98uswO962dhQUODluCDbpKE03MM27BXGJ248C/SWezDFNOcCPBB8i
Ti/uvCS9WagO4Q3SAEVnluhup2UI1+AULgG/V6Gr0rC8JJjKSIMeJHJFxB2qqzIqlS6dmR0B+FXs
B9lgOZ20TGXKrbo5tFbxAE/io7XFkWo0FTFtmPHvfJMJXYZ1eG2JaZe6+S6Nm/K7t7bI/HG1p5LB
oc3zVFMSBMWRJ5m8q4P4refyJrOe4K7UPZ+tpdVzsDuVrrI0dBKGqiFYZTtE/FOufJkeONORyo59
b0B+9gW42lMxxRNnif9oe1RsEKSetCK8fjcqg1WhlmTrBRLaxx9PvPg6ii98a4nhS8W4dKPzwgEw
+I6NtlIl9OxYxByB1gofVg5b4P+3PYduhrJRhO5h+g9nUnAYz967lcOUp+VxlXu32Dc4LLuzkb8O
zmJbrqWqi0vsuaga42D+Uo1Lbju4rEkWVU9UIHYKvAzbmu8MVCYR/kYHUbknwzJdgOp6y9iQoQzf
OuR1lwLSoPLyFJ8FNbiTS3T3bHomcWNtAoldPwdVO67aNnO4A3nBnf1A0N6IqtCrK5e8p2PjqYqu
lvSWfePkxH6H88ViA5Rw/ySJzNK2Djae1miO8LbZBEc6nVS/ZV/RRCG9F0c3sOW2EKvA3V75apTf
p+5QsztBVasAmNxrPnJXmK604hcQYW/6mKcmHdanlD1KzXcr4CDFpU+FMRziAJ75Xn2UOeobNfUo
kxKpf3xGg4lCbxR0nhraWZaGw8JkqBTAjBWJX0yRkHRibWFx+y27nN4Wx3S9aoZGE31vsWv55DvR
nA8JExtcgYZfK7B/FioFaVEEf2U7Bp5nm/Oe5hlIkeQRQCPSPX4TWljE6Ttp9oaWumLajAM5z1tk
zYqPDUXduWHDfQ47igfla3mWSMA8ExV9y0a00p+ECFp6iiWsra965p56wA/jmBr/WCsuWkHDhygi
IsqfBS+d0UkNukMTbRy/UwtyN+P3byDIAu+CUhPCtq5Mt4efOt6hqtFfhWYiHHnkVscWxN1laGut
jOlNDMXn9PKU+XN8iZsuwJNPBnTGp1Iadehp/g90eHTSfUFBCMdUfmV7oi0K3ExbtskALxQO5hJ/
kPjrvO/jkOGUbrEcHBrDUZ2SAn8SPp0Cr5w8r/HL4d92TyJ1+K6AG/4HIk5+2uGqG0H5ctm32+iY
ocI3aZATr15R59gaedvnyJIHcp8CvC83QODYD8TuMhnMGkl9dXPyHMBOxow4WYGbM4badRzy4t+e
DT8egxPyge+4UriZsrc+AXWtiZuvJKaaRo8WkhUHzacQ1AMOQnP/jYO7GdNRfc6RZEj2RjjeZPFb
BFo9ZCs5b3NzZ2kLkeYBPnYBtf6q2YVcxu6wLPrTRS6YpH1i2syn2/0ZhHN3T5Sg685tB84y4QLh
0ZG6nt3AHc3CvhfBqjwV71xQA5B+V5GcP3s1U4aWuwXPz9EhKEdky1mA7GBBSfs3k0Aa+8bn1C/F
8o1lYUcZN4faLHnOPDl9e9UwfBSShKzENkn/ezEuPaudkJDq5yCF1vNmOeUGXXg0crz1I1ZmL3iq
gEu3jObi/TcBpsJTY72rc8OC9w66dcltudp9ay8jR+9lCEEcYkZjaCCFvPxyEXvXFqql4gdDhrQa
yTDmcd8c9+33YHIBt+4p4ZlrpAuOcfzxI8iGaE5jv85whkHujX9sZVLZrFzvM29/+3PDeIPT0jD1
io5NxlFKjZvjvjUhJHxESGUBpD4RunfxnRJfZ0I+J2Bv6tTj+cFlnwzTmAhp8n50D4/EnT6okEfH
r6XbWduuZa7F0PGDmN/dlr5JSGlq7hyEPAp05mwjKcC3fde4T0az1gQquaqlqP+im7E/GlFD9ruQ
1PDp9boc0zl7DRGFOQSPLS1UAZjlwh0zyFBh0nLbnxADTl28hefcPc8nJUN0X7KT4RFwc5EFAyMk
q5czy4C5TCjj/d5wmqolbTmJaRXMRZvvfBywCqFQONf2+J5LNiE1VfDqhc7GJqrW4cppxXdWbTgg
ABhV4cleWmsH0qk+tLXAtxsRa5gZgyi+JqHN1RTwNFgPUBFtRRRCFqicQEKT7SB8AOm5PH+axJjl
zjQxHk1mvHxys/LR8XElxGKRkIPQ4f5icfRAr5xHbWVOdjwHw7v4W1AZvel1WYJHzTNGMPAcd3zt
MBkFnXU9g+6DN+Qcbj+Nn/8WO+N7a+O8l90oSrEUEj3mgP588pUaTHAleSK4lJZHZQ/jEUKZ9HrR
Ee0ybw71z752kWnw0mviOft5hwKol1JKUz/6nCwDQ1YJJVmCsmyMd0pn1QPvWH3ikkO45cYqA1sc
J0UcdktmvmncVZDxv/V8neTmUFnOzgvzB4TXLmqoiV+nQyCOe/qVffeEzIoJONPLxv/9VhPywUMY
0l/SjmFVyqFrT62MjujHKbJRG1dzvqTraD9HxLPXZ2cP1N4uCcU5FvewKPM2L7hELSSMZyA/iWce
/HxOJBDrz8Vy45q9aNyP45kJ9JmCmqc7VM/XkglD5a9HloF+2Ph5OSr1kK6J42qqKPk/jlyjNIba
4KivRokSHv6PGqGL8O1p+6oSRtrFwXik3tnL662eaV+fiavZmSfBYYg3w/V23ifQqaBB9OF7mfLH
jGrmQFHliEERwvdYDFjRR7HRTyVBELyc4HdLMV7DntKD3TVx9Og/Q2KgbzY6QpHHs8N17TOGQRba
jIJR9FjNNQqiD8sE3KXWXZsDjFP2rRbcPvRZrtfvEHBi3N5ZywGe4KbBhbxtDzwl08YPOfF6G9p4
deIt5ny1mToJsB6UiEEgzDw130pR9sLAR3VfbgWsFh/pSRC7B63zDK4EzSJ9wCwY1yE5saf7mwKk
0QOHowIgA+VBEhdM4cT1TMGoV/31xKcwuSJYOnR6DvyVZmtTFhdh+M+t1qkd6vZnjZwrmD6jBqA0
0IPGAD0LJTTF2Y77IEPZDtkPWrTIMe8Flb+cTLATNcBDIqDZMg2QTtvn7bFqt7n26mVJqoPMXi4p
erjUh8mmlS31MTCD/k/vKa8U66m+N8YkxJcRoQRJOEcNByswonk3Q5w76ckdPpSjA6LPYWLKiIZs
r4qVfHagFWt1N4qxOAa4qnortn8SNAbPM/zu2K1LPg2n9JLj2jXhc8CrnTvCUtOqlyL6fkjz++u4
XnhNKxTITm0sgwRpoDI4IpIJFjHkG6zt/ztqqXa3p2tP4IXBygDBbrrfCAFhqisr+swGxstD8coh
boSancagAT/xCbYF9qip7x3aBvSJ6q0o8qMH6zYsxNgjUaEL6M7DfmReiVgn9gEsex/xouqNRkdL
8mGFD1EC3CKLPK7TBXkyFjRdE+bfbfrZ8l7WrM80huPinnfPk6cng37yCPugnP8jOUv4oTx/UxRa
y/mojRDmczeUkmSM4MJpGoYWVICpVMSnq4xEOPTi+HMZ7MkM22niFFOIIkVe9NYuGbIB+KEvsLtx
/PJ6EsyzwMbL7xXxWKeVhUeKVwl42md5iJrUi5YcOQbkeMA1Mb8mcP4SpH5uNpVKLNfW9SuWIZWy
cnjL9rWJsDgD4ofVh1Oftm5nh6y9Y8fs/Qvl8vtm+V6UtPj3Aod2Xutml9h8FzVDfoKnCJRKb2hQ
lAAl52ETtq7n0u+l/75gVrQ5x/fOKTwAm0pOpcT/RnOAyBBOUpjWT0+e4uR0fQJgVR1swNkav31Z
J2HXPFX8DwBkgAkhTOporBBdPo86ixMKJKVYhOeYx9ru8euGhqOxH45bi8pP1ksfYtslwLKeVoUp
ja+o3YVajdcbjjCuC+9i0bXu45fT5n6u41nmgnpl3ofrI1bAePdfEkRAhYsW/iDnO/lvD3+XAhpP
frD+cB2z1mOhsQRBfh/iVZ4MlfSNh/G8brnWmeRSFOUXL0BGpYypqu5uDmYSnr58cj/W4f84BeNC
7FAf2WSW42HD7YjK4Plb19ezff1Ao4u38c4ZZPvdkYemjrcllmu0MyrQrMgBSw/YRmpd1mdT1uvf
Ltflk8rBz71Cd+XR1DKRFZShJviYTn9MWD8qI8ooqA1LoqHhzSzo3mWrwYLJ80TXZ+tKyVQ8koFj
ebu3VqdyXoc3NiUaQXzPgwHdvQZOBSej/oDezY6rE2Vry/9HgS/6KFJHEbxuUCk+Fa5E0hdrzChA
+3WYHQiUZfWya7WNWuXOpYF1Lm+qiGpwJQPd5ArcbTKLxszu2uF4t90xJ00ODeffPTB6SH+OTqPW
llfJlugVzXnZuImtylomttscrlJRPY2J8T3QgldvufoI+POdIfa/2RnJKzX0Zx0VUxiTrh64dfaf
KPVkNTRC+ylTUAVQTwPO8HfdhM+hT3krIgIXDZMrDy0JijKIgxea+wBhyj1EG37yiVYocAa2iftR
f8E5OrlSOlKtuLh8R6IOZwZMaCNsvMRRVT2nYiqalSWWwofHBAddC6Bm/HiTsb7cUwMyw5f+LH2R
4WBJyfx7WWUf+RnohOpJA5jxRyexpODOJUBpfr96AJrBsMvvAsVYNyTT5myWYIquU0YIgC4tmkAn
fEILoA8eSlpmVHmbAqlnmOT9qX4I7RyFPK1ls24aklrelV3aBs5WWXKCup+VZrt0SDL/ggUM8E/7
0C8LeR0lV+8hlcrSF4N/Pe6zGbhf0DZMxML26OLj6vz++pvUnBOwjXvfc/q/PJGlOgSBR37z3Asm
rhxH9sLXL2gkio/rxXiuEaZxTa4N3XardEDSy4944ZIOGegE8T9adNKBOUK1QOGzZnBS+YMpY+1e
Fyv2z/2Eb7A8TR39k9hocbjzuKCml6ls9oLSt2ER9xsF/RHfUd01deh7g1GsF1A0U8oa3uQ4aT2G
r28GKd0kqYK/kpuWbk3SaKaF9U1o1UUhfKiGTi00bEWKDlF0EgoVaICAYVcxl/lh7st/LOhtv8As
oSl6TZFw9r3ucf0AcoUn0dMYGHO2XQ+tQ6pQXXok7IcU27ffGr+L1W4Qje0v4khWgp5PrUAewHZ1
6ou6f5i9a76n6YFvusYfXZ94a8zLjr8H6nBQvdaFZ4hBChFo9RIyC0UQyMtoU7+M05ptDskCzDUa
dSthvYue2mUlGqvd5NRDKRjZcZssNU/KTAPQgh6/MF4neWN7CslNRoBvLEEZq6gfb8pA6DSmw1+7
8JXnneJoslzl3q5e/24+55wofqHEv58YHUSk3jJweeyWQt2HKWO5B+X/PuPgsmqYQg0oFiXc3hfm
t8mckhrFUPRTbeHijXyVeSGuXXFhtzSqCNTYqaV1++/8CG7iF8bo920cizWoCEoeEBCD4a3LjEki
nHo9hsD7XpxhwfZelakt4u2mitMOnQDpo3a6O9PQL8RmVd9ijkeqfQipDoWCB6e8kMzxdChM+uww
+3VpkB1QqzZ0t4bOnxIpst7PFsdIGloSRmFMno4uyxSpoLCEGz0Hdt2BUByGuWCiSHB87p5Z/O07
tMYpSCLN6+qwk8KY4aTuFCK5p2TajAwsNoyzioJVMVqT4/ZwzaUdpB00WUQQU6tUC5xv0KbO94R8
2i+3W5WE3tYh0+R/tH91RQjJkuGMyuKnRDtwc7kbTiZ4203o2fsZ1bx1J+6NrGugGq8+cPHc3i8E
GjLNuhV9++oXZGRC9BXRugDGEq8UP1dFx24bGGfi6i7y4b+wurOt6l8yaE9YeK4p4OLGKcwMDrOz
lEJ3FzdyDjght9G54QVRlVElnfKlCn/c7qE5dkdzeFWrjwgoCgTqGmrhC/tQySKp63wPzUs/GdeE
jqu4karVm8+TAfOzKAQ8K9WBoqmlQjz++uoU7GnCyd5mubFE/sIqn3g9c3vtDi3x5CkQ133rKSxq
X1d6XKZGv7fMEi37NSLXm9Ke2xaeZIthgc2RbFU2Heshc+GO23LQ5BFLzgUGY/FgL8eYVTggWUh0
a+zXboQezIj61r+l6S9hzxyXFmw0imORSBc3gijbwT3Y22pkdhlnXv4IEpw4BibIpmld/3U3ZdeY
gQtGmynCE39PkGDwM1fMvh8USkqLeTIbGHOJpOar28XqNahdphfe32zM4BjhBWZvwASPRze1f6St
rBdz8QPNVaeDAzGYnZ0X43HQxTjJ/3yYxKjsZu5tuu325xgf31fee1qckTomKad5jG/dnrgKKobs
1ATBsa8LUYtqaf+Yz1P+yL832MbHFYE6z85F1dRcB1PZLJQf4x7c1NTNBsOeW+rNieqoY8OjzqGS
2V3V4coTD71SQtXfCF7FewvYeLMhLX/w3K7woo2WcbTsbeNPoMaBbuQNhWUfER8AL4ug6fPzeo6Q
N4i6QDBKXODnef8pmgm/GwwAL4CAzieNIQLCJDwr+0pKtQPogOuVNq5fT5X9gEcvKtFhpAuIiTC7
TIuPEOPZBg1wiFIxXuu4O7UYhAF1fHShHHIInTr/LupHlHai3FIk098pTcGvL3B0qFPVJshSd3Vm
ivsPB377zaDcgsBhgmtwb8CPZKu+Ogfq2S12QAcqegqW7ry4iFnWP7V03Tcn9Ij0NFQDFnHDc7mj
5bCy0XOk2iRuBM2T7eQknmRCkyU8M7H9YMp++9BSCxZ57/PVTvwdODR96GEq31jtoY4Ip7MeGPsw
Bkh/MhTGK3DiWd7yYkVuGen132I0RF5cXvVI8/GLOeKCVbQ+aKiIfKZJ6tzOVoet9nivWIqqgFKN
UvcVrmjsjukjYWq/2G180uatbtg8miKyybmSFOSaNu+C2BwEeXNaKRVsZGltbEiEuGV5TmZ2Ylyc
o52oe2t69mzgWjNXksktcClb7sNLK7X9AWwO0tFrSUmREdlcg3/ph/ZZjKnaahRGjEhw+I0tH3Ar
b6A4ObWJDNkua/kjDF44nMaWCLIkVsnCO9S42wnrjCeVtdjyl4JuOSFJepKmckKv7sLmJE20Gd79
9l+rNvAeHw59nFairayfLZ1IGwqkDcU0S/vsN4Ey8BFcmcNAAKEkV0NCzJ6NdtOpSC4IbKHBpFEm
PZ4dGO86JrSFTLNySSkCGI8V1PdqYL5qdxTZB2nI3NQRjJ8cLfPMDCDfz91X+P5nJSsR25H/1ybZ
ZdHRC4ufeJqSDB6jDszs29RnaLWISOw/rzX1sqJjePApw8Z0hmMyp5DqkoKnf4ej4J9QEflZ3wJs
NOZ0n2XjOcwVcfNYPm81pmHOcW1IdK+joFhYiRQjXGXYENGPwvlHdb/8MSc+eM8JbYwwrhPM4n2s
c0GR3c9Gz9UtpCmmjDyMSH6DMClSRPJ2luNduxaAbZU7GY/fWwBksfW++Hj3bxILDg8NSSRHC7o/
VyAg6K9GmSRlgLmHdpvPGtZWzxFmfWBUl403RO48NvZysVgDymAUCWa4in79eit0/w9EEL7lI5Pg
6gGZJhxUWrE68sMpKYgdUPD1KorB84GYUZsb0o5zg6ZDekLGoGnPn25312ppzu8kurQbPFhiqdQ7
SrWKLsyD9PtPXZvGcdB6jbRYJ+PRSKR8WKKj0u9McsvpAUJztZ0tqdYD2bkz9SASSIulFgSh/r4I
umfLgJmLo1E2DJadvSr6LIpkDSSEu6sFfRPobXTn4q8zjPZE4Oxi2GeZOqFtRlMrJZK5JOGf35EL
5WVJGv0YPPbj4ZPob0BG+/tXR32JH4zG8agN7nRrmGIO8Ei9j3rF+Z0aOjsw4a4tE8pQneuqoFwT
WPiunQEbYAK2QZEdtJqVMNmPvPXZGOyIJVOpghDyrENDWK0Vu0Ovg/eSrPFBLnLXcmqRUfez3w3O
gGQRloLrKwBs/GJTCXBSAlr0ZGTXWX2HrVoXsqDSRZ7W53cyL2RRmJGQz1hhXkpJp5/LHRqv1or4
Tb/LrsJt+/4SeBQ+9ATUSkYz0T3KoTsXCoBdCYXIezCMc243rOUi+x0/7FAo0EQFX4QJR33ByHgO
zd3xPA6VS/3U6vCQ+o0SnLb+G9o/598JDUBLU0clHGjungErHGlEnVRo5xM8TVkjQBpisERonDbz
ODUNdutwVWhZXllAoALOVujtGr9AAnsz49W3p4ydlwFEDipqYWkYk8vBaSUurhpLnsfgfnS8Bpn7
tkq00CO0tta+M6XO1As5w67whefgB7csxp0SsE7WMRl+Ir3neZgJOVZpgKOswJCshmJpfG69PrRv
TLf1wEbd/B1oBaJ1n6fU/DYCjimhj7I8Xe4Hh6s9SlG615XIZLKzsbYEEvik1HRfvAeVh3gZoDZX
TnilWaYz/XL8GnGS4wL0dCFPWjdzbR34HCqawR3lSo4EoiYVG2NlSL8k71Z+fvFYiT7rnBHBYsoW
XXKE903b2shsl5jFFoMF/EhXHgXN8EeTtjw+jJKFUiWAWR7dJSp73T6RvuIeKYE8wSLn6U+MBJdy
zL5p8UDJHl690agSkYA0MJHMNMBVoNLybHBONTU+M4shR461KcQoVZw/XXq+h6aHBT0GoQTKPQbX
JvBvMT/S6p1Y5UMvtzh4XsQDS4qUB6VS+M5mKS2vvvokr8FPICYxtoEgeqaTyxRY3xQVPJAB3T3t
Ns7d8Y7c0AraMy1Xub9m5mbuvFrs+1E3h7r0QgixX7dxtfxmjW2zIFVpztSoTB2F2dSBKOJtO5FS
ztSBy49jiYsi5bXjD0Wv1AUXk7ZIkcQBh76ZEGPguSdazs6Z4UkNukSYVUXSm/fnGzZfBTD1lI4v
z7aGObsJWYSwLMiXV+D+X8qrSZKkYfzpP092LppSrUXpG/FbzOxmhPjVJYGKD7T+yqoBBRBiCy8/
qZGalJndo23d7SPjjCPiYNtAl7Zay7qZD34WYj60Te996cNEHAlgR//qeUMG/ES2amW04z1GBOyp
A5quQB7sFS/E5a2LIc/OS9jb9HEDLuDPOLt/HKlM1yPjVGp+UJuBM31P0G1ZEgiKrr5gFCNW2J7T
86USHNd9jEWhZZiOC1cyW8rOvbKsSwo/go/ra1PCSvWfn8+7LvtchCBgIwSxfr1r+2j2imKVVxS1
pkoEd6InaaWQ31k11/dL48F8CSgXK1uIT+196M5JFwV+8uYazFZU2/xdXh9QNGbFdmU37Dr9nkkT
vh3B19XozEoF7Y1OO9BfQyEJJxXVosWLj7LoufmjSUSIEx0mGoVqxCsSB6EVZVgj0sdxXv429wEP
LaxsJlz7en9i4pglzeriT+OfTDICiFRveZpqBbAAZxCPeNYN9bUoTGj9XOCoY6qzdln1JdDLD6wv
zIoMsb4CQAI8Azl2ln8w64rmpZc4oAIblcMo5GGGXYgiSCrMQ7nLcLeDUH9V+BovwuDMQsmuzaXZ
B0cMXHRflxjzDY8ftXVd7MrW+e8Qp2ic7GkYfjCvScDUplalFel30BHPMrbJxhjxfrXtd6Kq1sAI
tW1n8bdWCZkOiPaaFbgEw7Mnk7mpEqvI8SgDHR8JAq5pP7DQs9EYygHb+8BGRV4qmnR5FjUJOFbn
6vRxjbDStz0GiUMU8X8+QqawZOE3zw6+ERxmNls+zrp4FwazpJDz/LJYezY3flAesJ4Puzjx8HGb
si2H9HxvE+fHypRBrWPmn4dMjNHzmGy78T7xhui6gIiCoFe9E+4ACxb/QDF2P5xRdbMhTyh2R1rQ
kCieGmw1O3G7tuUl0IqE66oBX50BrUm8iQrXKrFLYZ5wxFvV1iqAbZbXj1j8qa6wfHTRXdr8xfSy
xB0DvQ6eHremy23p3y/Egpv804zh3s0KWk9CL3MnUrlqwevdviMa/QRICyLcRQAlqDi04KZ+zmGS
KhgSLBzvvb1BuAMmmBhCf1cJ4zRisYd0zI7yiD5awOke2dMNRZSVGce53SrlsinFpHV7S9rMvuXc
042aGv5Qb74MYmHBor3vO5oP80cWA+yGphLpZ46W1A6w4iyS1/73qhipnmmh4hyFWnguIWzxF2Q5
8gh4WR1AlsicNyg9x4/yL2Orqrv8xlk/UBaynGf7M0dkFwxsmh3zEsKpClfoxaY6N1WZdGy93JoH
JioFkY9rRXaRk11iDJlWKorfY3ANppK33x5vX/NdtWTtyk6glyGkRyxQoZDdk96dviYFLhCFZnQA
gV3gL8TUIkK+EdCRM6iceVYxSG4Xp9+aFkfw4Lt/C1rpcII0KCSR4nvxpPDoxA2qoq9kf8NGPHX5
EC1gpj4CPv7cSU0Ms7vzk8jGREWSau/KhS/SXWR0hbeCbGdr/yCto5dCgwOY7HltJs9tNGxXpITG
1+P1hxmgnDtYlVBInk0TpbKsAxRuPjxqXCdmmKSE8iTGv79SOxwxfqSBJJNs9HDKNX0cqMabpadW
SCOmnXUBMWcfDW3dldXZ8n5/kG+9KWWUboB4B+GlAnODQ9M0/CBBbwh0jZZNWlYLpTpADC4Xxuyb
rFLQuoT58Ght9BA9YxN+2QqdHjDWI7F3u4yWxxoBAZy+06osuleugOcCl08bT7TIq3lQZAJxoXYw
TNQWkiyF6J6tSQ0q6ktyuB4LDongM5ku02y654TCQBm+PkPB07B6ku4FYOJixi+nLe9xzeA3muuB
C4Q+UQUeeXBEplene0SiSuXCpmetybQ74DZNRmy6pY294omz2tgcX6imzgvEjpcKa8LCwGkizTkd
xNDNfUf3al5dsN4CZ6IW3YKHGR8Uax/cMiCmsiORlx1fFMJFRCSeC8dgzhTN6vbvzlUcVQKq5Wg7
V5dMg2pv2fMGkWryXIxfMXmu6odk0OWPtTD0DxitfTK3TYl57o9M86oPLtXmg7OE7znfPveIPWcw
Dh55I6vACqifMJyN5Jh8sFXPCI9Tm2QA8GCdyUbyGmh2fgDO+9tIVhCAqMXCwbJ6W0C/c+spD/SJ
Vl9IGhZEReP5vYACI3Mj+tlqOCcWrzP8ePh2W076YX032arrgEGbsRMx3G/6+YSA5M/pRa8ZREnZ
ES90dih9nHjmDUsjFwTh02bjs//+yBRjILoYubo41oKyGwx7HERKruL586gZxN/EX7+eXneSwMuy
GoPkkPv0kXANOd8sEVeCBWSSemHcRJ0urE1eM9CyIkPrrkQwyW96QTKO+6nHgJFwJXLx2NS5cG2I
Wq2LCcZ/DTT7lFIbOdTLvWNahD9oFKsVYU/RsyKyXtsl9UZREZGH7Bf/na0XVzHvdFnvnwTQniuU
pccCuRS/rDu4iAKUVJ5WeNdjHgiTTEs40UURr1sSi1yGHSCsF8pafIW73y+5PXXBP2cni/ZltTda
PdyqAoHG1uU3WOJbLOoo+3ttLPPIDs9jZq7EKXVvCtfUe5dkL1VtxIrz7JrXyci9TSfnQOmBgr4Z
2LwFNkH8YeyuOoioeHH//XOMWeHEiz2nu3sadTR30BgTiIoxF+yzHB57q3RoTIWeO1MuC5w9SOKu
uLo5COJTqt/ROetTEk14N9rEvBovun/DUTH7/yTXK+OzSYYLeQ8GhvceXqz/BIGXZs8DVqTQmFrT
ktnrpGq8WSp8zynfucNlzHWC5nO3spoX17j4JF3i1RiLOhxPBLqfQ98qwpyo4/g0k9SbPJWFIWS2
8cLckA5gJHdZh714bGv6fXgb0qKL3X+nRhYwm2V1EDmtJVt93E25eGhxSj2p0hSwvtksVI+1MWyr
SSqwVtVgapXsWFZ/lBaYYWZlzcHS7siCaj3SsP61RkQ7oKV8S3ogcaDyVTHFeiPPs4CTKWBEFrOu
3TCDct4aYFpSBdnt8JBr7ph7ofMcwqBIzhqiWJwO/bfohKXBS7JtqQVe+ZNb6T+yyrpQlLkxhpGo
5Looguw9XByyzRlBhg1vnqABcIRKeBskqNoq++jXu84WPIxwMUCu5jCFlOqjProDoXmyItqEZeDO
AnxRUt2jghl2hZYrAgrx1QsqZoukbWpRrO3mMxMMU0VBD6cWxmTGrGS/ZnaVOI+MGa9WqQNfrXHs
R956wSBUlufPy5P1c6V9XvzmjHjTFDKjSHH3JT4zMjA5baa/RXQpYUybK65kNA1JptQoapnI8RWx
Wk67JWqDLD9c6mblwFdD5BgwgjtihyMPaEte6LNCf3rvq9Sj+jr5QhM82biZOICTHGwKoeVHcd8m
1nGdNDKecdFFpE/F0HhhUMbejGks6AhUz6RMDYC6hg7gBVuDsCtu6aDbU3kSa3GhuSmLxo/Pqb0Q
OZBs1tg51koHC+lNMsqoRwKX1HKKJ/YKFOKyafm+Lm3aFFVRvDYfIMqRvLsWtt3Oh7qYcYjGlapz
lgf8VhLajFY2NKzGcv/ALrRoDYn+Qn5nabAX8zX8Dq5l4x2r7Wd1aQtc8/jVkeQKRJgoqID4KxFd
e4Dyzx7G6Jw8T5W89r1fUJ6FHCpyUY9vWCppkEM3gol5yt7WPjWuBlJgLGVwzEqeG+M8IGVlFb8X
8cIAyKyNMPyVBaLlloht2ThQHRcH9h3O7Uuub6kyPYFdWHPPqkaw4yE9dkQcgPd3BUmuQZNrl2ht
WGm+DolPyPG7rHL1l/T96GEUM4FqvACykzDdrFSHMuqdcBdG66RLhH7Co0L0RAfguieL4g7vcwqm
ZqwWejqBHNfPLof/PlgvaRbwxCvzRDBdgXX7ZnOPJ+7ZS08HkhdTzHxTuCe0e/37+rsoWEoPed5d
GBdvYZJ1uE1cZTtvdQyzbsGB+kP/IgJ7rMhh8WXKzTNFq9dql0D6p5QPXadLMK3xxk/yMElU0RMg
uYQm9a2fBbMdO5IOH7G5V+4dWWjN2qdxD6M7dw+bnJzBrqhnrBmXgqgv+EOVJryHl36Wtjd6BgUV
liLy9jbbMWfvpcfWfM0kQ0QQoI0GlvfKFMvBrqxi5ymnUBswcBvYQyTMv//LWc1XlyGEjdM40iKC
MpjFEbcgpijMwIxQA7tyd6OUaa2w7RXY17apcfyB9vED1UW+75ga/kdPCP2SRFaAdTVnvWwAjrge
bqDw3vL8OFSaLMsLvczNKMg5BAfyDHnrx8dk/33vU+RlqFlchs+avfZoIFsPKXx0UP23IdS7+K+g
J0mHD57iRGOoTM5E9nSDQyq954bzztDDlpfVRFgtaroA/YioRF9SKlkURZFR7meHfbxJW5wIxLTA
k553PGIXUkNOd8BQxLl9OTnIFTFPdkeU4WMJs3z4356dfM+tq24XQevBvaUcQ5GbWLXVDOI0GMTm
qUjoiSxkts4y1GGsa3EaCaBzNStuEYupJ+ClZO/qNWFmoH8BebJrsxAkNBb7AszdyhT0LNwk+bhX
LPaw8pz+x9Z0THOtwqJiFZIxVY8EBwtr2VYFGXVYLtOxkngGGBfEb5eUNUtbzQFF8FHLpGd96xYM
9e/8K0lMNd7t3TG/yE3Fsa6Ee4T73lA3IOtshzUewSee5rcZvbc/MJSblFzDY1usrkV9/m164FhT
tt+jOjQQK3QXiTSxpgglFC9vUIjETSipFdlHrowZLOEtyrko4ymGhxTSx/o9rBaGJgaFOeu9Tqg8
J9gBruOYH0LDzsb0flzKJ0mb73wk6Cb+byrIFWXSlMNXL8wq02aLoki4mCHgJWF8v5MYHjjGBEA3
BTa5rQuHYtKD6essoZuEFSSGqiawtzy0foxJHagsibEBrscH1emiP8inQWdxdSoPVTg8xT1LpubB
Tft6ge4KQQamQJ5jXs2tKCAjORa2gKNYWdz7W3PS763i4eIICiwLpDDn2MgV0GXschF2IvUNOxMQ
8TC7qqU8YKsuHx92i2yYUYnt8mj9ZRhUDh+cB7uRWBH0WY+h6h7kIWVeXZIYEIkC3jHt7gUZdMgi
DHWPMcb+bb/zIcvakh8BdQYZMlNnK3kBpZTe8k/zph+pQRjoRCRj7U8MvRQz5PvRK6d+g/MhMF+J
hhxdhKveopVSk9aB5LxzdWkKD5um2l+xZJUStTlTzXuvlgAHSDgwbU8tue1aqYTooMs+bgNG0soT
DadpjpdOJbrSuR3RFcKpiok1ylJP6gEt0WZvGOWM7VGDNPPYC05rXyWXxUEj1ud8vKZr0wZv+llb
n3wJXw85bOTr/xukq48pZMTqNvZ7hgpr8X8sYEQ+19ISHhYQKM8UDR5N5hdxFt4WMeJ0xq/d2w8J
fGFqOSKsLBJTAqknlJSk8pvluxJYz6M07qQtV3pl7sjVMc/+CHbaEoGfkbJ3ud6yCprdgfDX0nPO
kKPuIT6hMv56EAFPg3A964YmVpiTJbjgSRLzONdCh5yjT7ZXvsftb5E+wR8c7K8YBCfnHV3gfXLw
o0mR4H+s3Wp6WgjCz8FmNXSM8isVUx/BU+5yMDW3aKv01EHStnSk8ckViBzizqa7pDn6BXiwJJe+
UjGlL6j8vxUrvJve3X078+z37NK3h11BmIApSAhlwd2eANQa6nrw/NipDsWQ55t9JtDj3Klwn331
lDvop0LgbyIr+s1IKxoJEG/NOKinFLgQfXN290n3UzXtyuigAUfP1ltbj9ZQWsajT8UO9J/URUEj
6PgtlJMylqDZgJ3Xjv7KdYUwF5CG+lDmSDRC5NZdxIRcs09o658UB54WdRRrsi1HCLLphpKwn2VJ
zmVrWZ1ccMjSUmmjhW6sCL7ow29buEpGPFlDl90CU6sYeQVSPhlny6ihborUNUKbmNriZoLrT/v7
ZXXJZNocjfzJXIwiWmsyepjuyq4A4ugyYwl+tLXTVIeLAsKj4txGmhgDl1iRrFL4pr6cFYITp3Ok
liGVLtOPcTxysEzlW7OBYgPRR4+j/+/HERh1q8P6S3ChS2SmKA33Qg8fCBZNFlUojE1DXX9zcYWw
xaqwYLKQTpM1csgIYOnxMTcSl7fLxg/xz1xjVM2XLnwHIoIPJhiq3yPb9d6fLljNAgHdiWMEvMC0
9bOJyz1mLdmm6xYOiCYmPCNMC4GRYytwtEFFOuQW5m/SsiQ+SEiH1K0Bm/NnKvCy/XPHOkuFAe+4
QoPPvCP2zgO1xQhLSFqfLz84KwGaSHERqEqiGcgmLDyIJOPzQOQ7CoOk0/OgXcn3qwCoO2//j7E0
WThaWnWpw080NZ1RElz2OaDXVFhj9S1P/1Y5Xm7bTxOfeOtssts6BSK6zSJXitxUzahD+l+YO7OI
gOOOYIEy/ALy5LOvIp6Enoyk4ft9fY5fy7Eqw3gJP99Wg9+Kk+w0OeE78Il9XZroTVO1YmJFc9iJ
5+btXJp/arVFbMZFLS+LNbSzH40JiiN8rqCHggNhdokMmxdgqDEESorc7Gnch1Zifi8l/TFVs8tl
YfDKDAtnAFHt6NsPEQhR4frB4MZNpxoX0G2PLjrTxPxC4bv8fgNU+7fwB4qS1SnjGwrDEHVvXlTF
Pk+LfeIBelZ56OrwKtb8wOfbxmouezLTmUDifhSaAGnYj7vIdJWBKh+TAVwSt4tHNskCvprI2IYQ
qN2RgJPKxMFn+nxLzYgMncKFJXl5+0amEKzZi1GfF9lVZ637eaASmagSFyFuk6iMi3R0TZk2L03c
KPS3k+Rm9KyOFXYDAI00FumlvdhNm5NRbI2Q+NRmxhzen0AgkJ2++ZWhdIRNpjjLVAkaCB3m9LVc
GE5l5F4l3WRrFaDHyGeYVQh6EbFLkR08pxmDdpcf6lH8zTc4vJNkJwDrMt0I+QZGjxlQE2DGlEEF
2BGcMQ8q5XUyJ1cvHRmCjiYfNlIPWK8USotsx2RIFrVv8rnauEr3oR4L+gLLCEJQWchps8RTYgU4
T3tf5s4c7jnHDIW+4ptgkrs/vyY5DAoQZgfsZ+b1eEb3Isj4MT+wNxkTA61I9k1ocLvYkYYmuGSk
rS2mmpRnN31BvfXW8BGyRsCucxXHpCqi4dDDbraa50VijiFtjEgFOCoCbZO5KWc9kjkdFkL3juHn
FPOxR+TQlT1mJaLHgS18VKouDg6wCE3Ki2kfl9iX4HmShem9htE805NUWSm5lJeZYoTMvfH8uQCW
noDI2rWHkcytRBigVwtj/SSWaLdxTn9UEqou0lep/thyHnnCncKTicWyN0GCyah9E7AP6UeI+pTT
7agoHd3utk08KGi777jkuylANjVrbDBWnFjZdQ7SbfRikJUd7LWUd0sop1v7Pa56xPmM+D6BVsLS
1VsVPbckA3j2/sKPfn+FjeyBZyYQsGUK3fbbY52RpJ31ep2jjbTmnztfmFbJGhVqAGv/A01XEG7K
xEzH80oSp1sITP9iqkPytXv/QiUegb9VgMT1m5iDGMi6rm1DLaNXr1afPe1VMcTTQvkRePnsB+xT
zM85yq9Wk74TfKDcw4GalqGO1r9XbdfhU6iGsqcPHHArWg/VqHiFNIsO7soK2+4wFvJS8348FmDg
+Ov076k7yB/Piw7yh2CuR+JInIKI/O/x+NKOvQu2kd6wJ/X32c9YZWTyMNvSs9ua3X+f3IrT3KrO
eFf9taaU04rHbQUzyd8ZrLbYxsSH6BeViI/3oZyFwmDBWxpW8iQcj0u5gIcKKb3R155BpNZvSsSZ
wLKtXlTftcsJX4OEi+U5Y8e86Za5DH0Qot6h2UwX6GCqY/lq9h0FRFF3ALYhkKHaDHDsRiq/iZq+
6ymuW40dZcP01cVSEkanzZwcTMwdMg1C+D47PB3U6OmLHUH2EwC7C7SX4r2SK/B3m7uLyLP3vZcy
RwhL262UD2T3SecaJlTtye9wzcVe8wnJJAtsApQqd1JGY1CtaavXlvVrbqrKmRYtbDegzkO5ZiDm
VLyrKgWwPH2VAOwrZU0tiVEtqgMyZhTPx6tcQhZtDYgI2+BooTnbdmEBPjARQKV4gOlYAqUqMxsc
N0zHu7u0/OJt0c2o3mmJANlCEG9a4yvqz8y9H1f1lxrxfXCj7jw0iIlt0c29RAdOQZIYkkDQfxOX
g24LV7o4e4laiLrWjqUsoU/rq7SrMqRKtf6VmuKAlAfSlAlE1FhieobUVl6ofE4L9ReHRC1NQeE8
Vct51bz+qFuSYTvajk2xRIH+26hBAkkm3fFK6Pv5k+QPZOQmDD8Lfg5oe+XwHFuezRZURIhpGvky
HnmfUtU2TAuObY66V7ZzWEn4hzCBAHOgwodgARWQkedY1auXXkkIYe/p2k7jzxZ9os4zAg1L/CIm
nYD1OMMjTh+hFPrGgMWVkwhHUvxxqdPZ0u3WRpjz7Z7rswnxVLQfWg5UP5/3Alc+VwJlsM2p3xck
xG3GxnAXMhysRBkJl989Wfr2mkXty+ypWnOrzieMvYTSPozLU0n9Yo52Sd1IPLDhpf/HXFRjx11r
v/E/V5Nyk3lMjI/9KmI1YrA80O1ew5yIilqxA4z9oXAzhcIdtJnPdGekeqiYSrS0rHo/siQ4lLHs
9EgAyMsrqySrTz4Mlmp5rzRBMpRfsEcqGwhL6jgG3UVVYvcHHy1Yzv2tJ6BJwmHzGG14Ip9tFEQ3
ld2xC823LPGuYQCs7ysEKVMuipIC/GiYvYdva12Xul0Uq3g+kyQ97KEufOjlH2gjtIPvcMs/OP79
IOryErMSF2ewE6C3MvNm5wzH2y3mhnq2scPbWq+/T+O/vDNEAEonID5/f0mYf8z/e4bLFDRLOvN4
BMbJfzGkIvMey9U8s0ISJvp5lKJ5w7LLiBespfGvh7OBxERMhkDaUxzBcoaLL9lIoVmAu030cUnK
sb9LayqqTeUb2UWKyE6MEW2q46Q1K+tKHA6xWY45jbQSOW0RB0v3H65Qo9fx1pheD9K4FOEXme9X
+YJ9iwBtsw3zwriMKhBnMxk4cclk9QKsKy9akGEALxxMmnNp2JAaVcnsAtOltn3vall3XE+yhCX8
ecWaTcEEGp/pfmB5Of5Xy9xxSD6nS7aD7n2h5NhT9Hb4CCxOjKlZnLOIVAVZjDaUPyJjZN3ORiXj
j5Bh6zusq+YqlqjXdhUI36A8NvPqpRUqwSF4vIXIAWnbMYZgCLnSjrqa2sb+F3iv8t1dgq+9Z/m6
VmHdgHhH0G48wYAeN/nxGHv1st4iHi1BnsZMja8VFOUdzDjc8MWcohi4UPpZm4LItlPC2oUhT5g9
nUobXetrSLuxKBSLItTg0Vl/es/KiCoJ/t9QW0Y1K8uJxAhnjea2Y0I0wGYgeL72YIURSe+wfEdl
an4xoX81FG9PDJosicm+oCo6sQ+sKUI8QAmnjetGMqzakUn0iBjpcd97bmqbNZKvKfuTgAHD9yEB
W9QyTbENm+DkDw35XvT7wwXM9qElYqmPqgyDq8Vrz9DpJpUxlhh+TY2TQFqpdmgXRoG0bBFfrU0n
68mKgpJb75c6eVtBNzAys71zUNTxI8jyI9/ZgSgGIxE18Nv2qFjJNiXcJW8iujOX5ayYbnRoV/q5
+ljvC/POCsHsXuw9p4pd8yvt+v4v7D7gobD8TQaqu0W4WHWBs1ZwFnZjaPYZpVdsJEmKUxpn3Rpb
XoibQGyvqhV/c6/bAx3+dIH902vr2O8j+K6Y2dYPxCPb36be2CZofwnlAQHaIY6EPUXqP2BrS+2Z
CbZYAlQxVyy6JsW0mXK5LVbU8OVy5FxPC+nD5BBx5QkWxtxuQ8bsBkhJSDrqA+ffnPT8hzaASiiV
wHBmeVXoBq+Ux5J2UTN359EiPkTF0YVVs+oaCeEdn+6BqyhSbE0o7ArrL6pNtAPtKr2Aj9dhwM3A
6+DpPH/yOqoACEp/P/8hxeJgEBc7Lw9CfRWqIGbqdCcjDR3Tgy1VEDQ+JVseIk93SxWmMp8QzUV3
oRZOjUdVm99tlrouMfqQd8wxQzXfF4Pfzp78lzNJ0yjN9mGj+PmBB8ylpZP1BYueuvDPDw/kLuu/
3pFzFiy16pRqRbHEDn0SYYJszlu1aKwje4z2ZNBsGbbKTZVOKi3S/4t5hb57vjeHiq9CUtHZ4j4h
tpmZzi70w9U3gNGrMbXTSQ0MQYmbkhbWhYlHpNb09WZe1rdRKDM+QZ7M6UdvNxaOK6bmdooHS5Z0
C63RGEQDuxeDWnjtS6vL0Sqe3JnZL3pIjQMM8cnv8NG4fCMq793fl6StFurHP4k8l9HaQuiOZ1tB
CjfRSD/MnGtlIE6NqjVpVeOMb2Ku0eRqJb45y8dk1IU8KnVnabz1bD55fQR6Oi2ns2jC6lZe9Rg3
RYBi/iulLFMbKRGh39ea9qvkXB3px9KZ6lWGIORpYsmu/6ShO6M58T8xBJiKquL2Hh34KDNomvYk
67Dt9UrwUjYS66H0AqnS5d/dkR1A+ijDkdvq8AUHKo+CqnIipS9Bu+xl4qQudscZE2djXm5bcYfM
jJymQSgSO+Qq2LGKKu5uJmBMRJ8lZIaCuWX5Qh+xtdVTtupfl3L8UZoqEZ/LZ65SXQJLYdKd3btp
Sg6n8iQRBigznE6gdoWorVT2ds/qIeBDXoPhOf6nFMpd5cCwqZdj3IH67g2udQXDOUhMtPxDqFGw
UcSOuff2+SJLTQk45BhCYL1zTDQdHZdeMWkkbCSUjo+n0eq+gRvl2a+usx7jYNBTnBSS/buoVpiM
xAmePCxYBAw4PJOwvkeNavU4fT2upezdQD+JYT/jDey/wJEIOvh/aBkB5dn13EdaZF0pUFfSmblT
xiTFcX+n+iojMDFSjDTZ8KrXi9UN90Bj5DnL6BcPo5lEMhfhWH8otblNy1ueGiW4xifWMadePzok
92hoOlvBDl5Tlok2LTCbnBO/3/eslWkABbyBZcdQ4nY5Qlmt0VFwqwe5FrM8l/RriYNK/6HgwePm
AqJteEGJY1s5pSbf/8M49+koosOLhJYryrE5zfC5bUKcn4QeCEBrqVVBFKZ/qiP1Xpo3bWhWELlJ
lQFpPkuocN8I+7S+xUk8V6VZLd+yAi+dF3djx1toKWpbOiBPF9SEuBZe1F9/W6xFFVjVTAfySVF0
Y51fySL/71ndU1UVWQVCZR5etZwKuzjpHN9Kr5LrIHAXzl4T8TqpDp/Aaju6nyMeY95zez1zJwcg
AXm3P0E8sNIiuzFrAVQ1Jqd3PRSh/khraP1mfHvOlJtF1stfx98N69yPxrz+xMsmD3enkrOGoHz3
Wz3U1YTDrDlLhjGINXJMLfIMZHdWD8pDRLc6EctdU3xn0eV+34RtH4Mtm+fOEH+o4zIjPSMh3RKA
NFT9f4hTZvI1vVDoZKHRXAeYlcZs+OEq/a0azKmDYjIdOirSHC9G7vvIuheUh5+24huxURZVJfLu
k7aKyerIf1tkNinknEg6iMcndmgt4ppgaxdjFkmPzMamxvA6fpegPgLOX8GWLAQY1puq6Tptusp2
IxmwZNLeAn3BcidVjhVVtnKidxUELh3D9pr94kTVxXF4Wyb5NvfmfIRK7NNtAwBq5xbSf4t8+Wlv
cfNZBUaWDVPt33PRpnCE05tDdmRhjj/osNIEAWsJe0+c8fTQb/p85ixRW55lFklTYeY9ntQhpUUM
XJ4VSr+Q1PZNLjaxZTKXTdficj4WtxnNexv1sW/IYyyMLU2IvsP4mXM9DaxHoS8edrbu5Ul+Pkw3
6hicQYUQsxDDhMr04ce6bhQOAeCGIQ1zt6EpNZK8MNslkvrQ2JxkdLOLrcW03KJsNbyYdHlqyljg
ClomN78SMBlmoN0z7TeMxBsBgBoUIdz+A8TNsFlH6P7ZJhkTcKdgM78uSmtyPuOQPjCvkPiv9iqm
a5ySeFWBHPjwF0sRVGgfWT15nSDGl6HZw8D/b4Smys6RVnDGzOZa+uRJF9FUIY97qmq6HuJk3fzH
xnGFL4oPySiJZ3ad/b7oy/ca+sniZfp5yNq1X9oUt6ORy72Xar7rQ+92bD7hHjLBeJSr5GT41apq
ECDMgm70zE1UrRuDWflnae3CtF0k0algp3WEBXkPQqe2uQhjT1XaLQhBb9Ye5GFeC50VanFI/G6M
oHjRqqnWobKEbxyhB492hQStz3K0FZpU97AVwtbr1ieu/Jz9d5Emz1EagPmt6XMKufcK2iOv8u0q
5lOQBUqc7nDTfJTtjuXqzp5ApngakhiiiCbt3iEoRh6lYdqm4gIKZHqVruf9kt1+XwGn9Aw0oJYw
aOJYKWpalstihR5xiRkciRQUBbGQext7Ukr3Xb5ljWV7M9gEZAMbWdbs8rFI6z1uAHGES6m12EHT
AS6Q08QHyF1oI9JcmTX6o5vah1zHLhUu2iyDzQrZJjDRHyJ+bZziqduc75sEK9tcSKuNTiPo6J2p
cD4CnGekW/dxa6SD7rflb5q6VmVAsubdobkHfUQvU5cguq3d4c6e8U+G8cAOwIGXnS5knmZC9E/6
9k8RJoRkeZmbZrwVRWnrAfBjG9Tr4kLz/5Dcc8q2nQdXkXlY5jPna2BMO7icRVY20NeLOVnNbPDF
+PYwgzV1yMggtXwYBrohTsDRNpHvygKfunf/AmKGl2d+PZfx8xIGKCaDxIjEq9vsVQ/sRcsvdd0n
YzRigB40wv46NJSdNVlCgoLtN/LF9KqvAajZt0uPBsB6m2RFA4kD6aHYVZRU47BJSYc9VSCoF1oQ
udDg216/xBALVoxwbLbF050QjIV0eMY2VmETmyeSZZk+43CBnCs2bsQQiRdsWHN2QYgF0HdqX1jk
eRxEVG8luDKtoLHcdrn6s9w90RV1e8RT1u3HA20zWi4V9+nQJwICLsonIL8FBxyLaanzWYIrpJNw
QfAkqw4HOlkplM1xTVP+qRC6mI6jQJJ+1vf/ehLt0x22ImhLb+qPHIWQwnYh7LerSPbk0sOoX0ks
by0GvDtBBlzAVt7C3XwqOWoibAD7GNzEHmFbJLXpC+Wwod4I0Tnm9sOaweh41J2g1ulIj/5KmwBc
meWsz4I5UmujxKnVUrAMsTwi8k5FykqwVhQff14CKev1lyQ2kBHPDksD4/CbgsPfhv8f2Hpgg58m
1/od6++nrA5rZTqWA5E8Xvd0FDDadaT65uj8rdTLRbtBTOv+DHWx7gyYsS78Re61lCbsC2QHqs/t
FcLYdRhJeHYb5ZJHdkWfDTImkv/wlKLLgKlT7Oas/Slc2yakAf/yvHUGGtdic6Rs23zLA8azeazq
7OSH6I4cS5PRx5c8xW1snlGhWUb+Rjhk6n/bAqenxam/QTB9znBYHoPjtst29POn8pi3RQudCkla
Z9c/8jKHpUTAuVS42K70BeV+GDXFhXyQLc4AotEkA+w2j73ISw/LU1hrSu9DgPoxUkyGugZIQP4k
lP2RXRIU0mbpTmZboZLDl4ISThzhKdRnKUAbQOX/aZ2fvq35lGKUfw/GDvNiWBxMgxsOylFKOwWM
lsqoaROv1Ca7/ebKpZeVYkNvaLg4gdJk8lyDlWtLvVbz4RyK8bpOY72BX08UOXrJ0z+uc6aU54Yi
ejKEFDRL6QNsAJWQ3k24WnC0Jd8VeEeiL51i2rCqKyfY/zbpevUwUZHuFpRZQZMa2q2642wbjf8s
ESK8kmTk4AMLqKRsOwewrXHoJyFm++6Pj9UPHNXbk1QHWiGGRHNIQNhUjT+XUZENWHJL6IswOHGU
PVsEdxmnS6DaaZnlxrJimPLr86NlaPeZYbmrM4gpOwL3b1k4XfLwcFwI4fFm41Q5SKiT5RRJUtT3
UVGpufFj3ShO/8SkVWzYq37hOTZ0SbMSdW+Sc8RoJOl8i7vLXsVs5boQyXKmamxEPSHoLRzvOJJP
JLloGyY0byTYcZLm2zbVYd7WVvChA0WOWm11l+KYs1j6axbtZGhL6lNSIjpEaaPMLhTnNJJALPDc
I4upTtFuUYQMwOImF5H1G3Fg4oD2SPL1p0JHnItgXsF6iR4a4QYsoa5C5qayOyeXX9tV92J2jDUk
S7YuaLUWnmql9FAJPvIykQjECeLYs0QsdMZzYLsj8JIIsvWpOsY0dgAOH2rWG4D8sFKsfk+h4JqN
S3rWGstJXc9OOtJ1ukhBmyZu5RB9QfFq5J7BrWK2qgDsndUxd09ofpBNM1V/WNhOmDWdso9dw0Kj
8ydxz7cprheMdPN8g52TYPlm+Tn9vLeJUKCb2oWx71S6Dlo79H+Chq4i8jYf/k8+gJHfJ3WsDREt
+j+b9vGwcNgR7E111fwY52xfKWIb1p8cCy6+IjiUaEWo5HLj6du4o49JbKXNek4CVtolyKjdp42v
vJ+ounl3Ro6mjVdvQLjDz0XQHBu/kGzhQ5ze4dbWXtf4pKXZqUVYR7GbLILXOxxwK6OoYZppokLI
UVaNgGWhU7DF/2JrZNBbkipDxMbwam7ZKuPe7PDfyCfqMeKfTJ+4VbxilB2+/GHTMAwsUaBmGd6t
bcuIuvBUZlCS/kwF8Squ3wxmF1mFvqXnn0Fjd1ydYBBgH/igoJytxg0Df/ztBN5mmeHbBXf52C77
mBg6xIIZ6qTRY08U2UvcS+TRtOCOqRWl71WJYQzHWeTchvVBncUNw6UEOoi2GeAnGgnkexDUCRZN
KnIY5ltK2813smmpKl4U/eJKBFe38nmFXlD0i5Sv4P7NbkUDkHJI0TKq3G1dXcDii/0QOrwj3oEk
JXysI7ZN7kMIn/AcncTmxejzrMgrvsTQi/Yvch7TodIBCkSdEvsTlSjP4J46//lJ8rTuqz7bS92v
EL5IyJ3xXMvm6FpscA44/bT34eTPAqee11wVoy2W3Ql2nrmhVe6B35nv1Kq59DUppyKLYXBAzZhB
idELn9mCjwb844lopgiQsLNHN8dx8SNlMLLRn7iBXGTqUHXfCoVhjgsmbxg6XzTHaL0dP2gRX6OQ
D61SnFOkxBSHcec1hOnDRee2gSu3Lq63gVVyZRlzM7+Ylty2PCloJ3u61d0E47hQASTKoUrAgEoF
XB5e6ztlmfJwfbUOADy0l8DWJhFLco38zw6rC3bEMB5waqOLeY+YUQd8SuV28rXhqtf4YIuj8Fz0
viFRVWZUCmEvMgQEXkS9+kfBf9yEMELKc6tODyo6NTQimLS1QrIfREZp4H4OhiUefG/OJ4L1Otv+
Elc3jbe2e2pCgUsXgPgLjFkPe4+Eu9WgIZXmROLW3jfvTFjkxv1x5tZFAZtY/hE8EG2JsZdLmKTU
r2Htwfr7Tgt/LofS2qbflib0QylqW5U9Y3ileQo3iTtgY1dIoU9JJgRG33ueNfXVEbuhiZ3d7C/+
gNKuRv4RQwwpWVNTqh7IZJkAaApzPb9GpuA8EfGLnn4hjxmARf6Pbx6HS3VSH3+HCQvhQgjF9OKJ
aWgJ9qbHw9g/cH9d2/CpvkDFLzqKtHW2Gu8oj87N0L7O4B63trYz9ry2rOGEXvQ7tx6Y3SgpkEdD
gcZSuPE5i6zm3MIcS7KCgATkVKzka/8DcqQMPMZWxqwp++ZMtJk4kSVB5jK1pATTIQLTYIQiPJiV
zMBEIWXWK/npGnTAcYxCYLmAExVnJl23yS0adSd1L3FgkZWJ28ed4+f4f5cP0ue4Kajt/aIS1ZVB
PhY1ztABlawkUNrv5DqsNw2YquLRnzKQTfI32QZQyJPuvUV1txPFlvE6cBpI4Kb4akPOTdUTwLzw
OPlW0eKlZjc5pw9w+ylYWI8hvw2I6MkLwJ4hiKJI2C2Mp2w3dTYAt6+TEgLvZBo1HffiGalbKGjt
rJ4tYHnYxFZT7lpz5LKL7f/StYmFj/dbvrXPMuLrAJyPG1QYrMo5tAazoY0oRThMjC1nF6fBGMZM
ufiiwj3jXx2PoBGzXugHrBzg4GE0SU+joU/9jXSLa+spBW+Oki1bcqQIr0yUs4/+Brlu1vpiZdW3
MX54xaMlse4S0gsW3Q9lFhYjA9rY21ZIdrRHM/oXSR1UJ+ZOGBTOd4DbjsCxegoQKeIY0qRXhUTY
y94IwryaJuYMKw0HxEF5sxWNAXY/c+xDcySPeABeXvOL90mFEwi1wQNwiFuHBDOwWQVdfi+39AC9
2mlYQdBOig8+JkqcvlNTmjJW/i8bjx5jLe0F4oqu5DfgNzV4Bzj9bawiKKEd/DfT5IcVhpMecsZo
36G+euVJoXEq4VuV38cPvSpDqVQ60IdyVzDXpimV8VGaBn5rS1MliBfys2IkdYkfM076GvpPauDs
7zcttmnqlyZf+/HfDXqG0H7OvdiWaEfGWfLXgN2ivZMZkQWbyj7rf5sFWTpbUVaVJHQYXCBtTibY
O8Dp9Ik7OFAeBFcS4lb8Bwn3hHm/icihZE0eIxtKf7s49w0ebDCqwP3Y/uAPnhcKdWkzVu4Jl4/+
krECX3Rf4WJollwXkbGckdRhSwGOwSEjYnn0jxCMj24FeV2hINQc5TFCY45oSLngunudJYT1qZlu
q1jhAlkzhrfpxUwS5FS2FrdyD6lfVTrE4Zc9qSkKucVUTyjEQQoR6HqxP5urzv6w6L1pNRlQWDED
zs0KdSXRvez4SS+Wdgh6wougpRrAFeRZF++oPOyCfIqISLWdXyU9XWCrAHHj0WWFpRGv/jWLqYtI
prl/zMhwpHY7nizj2m3S+xainyca379Tu6I2IuTrEhDfyUdU01edMqKntCQTSjo7pBR0dGACtv2r
ahTm8mzLZ9OYMgw/hnJif5Wf56Fuw8hs+B4lbKMCvwzYa5tT8AES4lfkVTa4KI7HaO2BDXruh73f
8dq1w7i76TqGure5Mf3gK6B2T7kdCVTpvWk11YVXUe8ADRec6nCdnsq6SaJUHlvQyg3y7Jf0cxut
1IXrmhG9T1WJxqV8SWvjKu4RZ5XaEEVkgj7Zme0dk0hJn2EkZVvyo9NQaWZfmDxxjYmaOHZtDTod
I3hxLzLoX/MSwHrNeec938XH+798cLj05012qh5bTUgsn+FR9ZK6Lq4zjzp0+A9pUOE0Hwo9ctDS
QoHVyMN/D4yDPwEPgAExbOULbrbHAxWok00qW0+hcIBiLjWF+zzsv97XmKo4WdTwmPHdOu6Asay3
OL05Xx5a91V8NBHl69renLXUuQMl3ugNlzb69ust1aZy44a3vzPeXnQLO+svKwKqMKLu1nvNo+Xj
oSua+Q04seor8OydN6Okr4QVNh78gS9AU27SaGHBzAqO0YurrWTrvFxIl3ITcsTDOJsn3ctjG0ad
6rsaSKhN5IUa2K7vro7Y7UvP6MpiNh9pCQYxYkkQlC09MhaLhUGVZS9DYpmKGxvBoakUOERyErq3
GJjpGcUcisHJs1HdaT/TXS2RQp0zA6O94jnI6Rdv+dsOGpQQPYOrJPZigjrxKTIGgBkLPj0KXaRO
AZWMPSqUX7nFFJRv/X+FQD4rBikVQXiEi5PMq3KeTp1b6XnagPMaZVF+LtZ7uuxkY14spv6Fj7b4
hPg+gpvtEWAbtj7qOlv/rAQ1MYSkJMXslDv+5MyOtzPvarhTycBOxjunnOGDkXDyHlgLLhbs5XhP
RKKDd9Nn2pLebeilORRWv6Bf27eExjn1Bdza2WcGoS+EWIlWaTKwvf4I1ijqSwXWY7E6jphCtvdj
Npu1WAyA/2Ag8rzCJpwvRJa5EXHwl36lvzyLRKuJS5Irutp6dv4XLmAYH46uu9i00dtub/akQl1l
DhhUiKEL4fhVQu5alnUGo0Wohi2SHn5miPfb9WJwlqr3BI/IWn6to0CJ6vhOovMUpOVsjOHcYbui
lmqU57tJFurxyMXMNmoUwjVmKlm6Zy7lRzrT82yVyWkFBI/+HgRF9T6jJVw6b48RU4qSHP7gdN9H
pEgZGgBwSLPnLGGX8uIuAtqIz2V4RwtpX0IwzT/bGa441yV+T7eg0oAUqgwCjMK8dmUvR1aWD7/i
aM+IVxEuHSuRsH6qFxoATgLGZNQd+5OnxFI4p0qOaLa5jEKyog3JnLfci9RxmDvmJlXZ2ANZIlbI
OmI50Rmnx6RgwwVbRAo/nkJ3QRGqslCmY2b5Fn7pBV3usFjIYJ2CWe9c8Jr0XWBwJoOuK4/TTT6t
rpDa8eTEz7gnniYy0qyZpL2qP5jBosFdbsp+CbHAQ0jFG3y9KLDlnVLteq8eAgaJEFTCa2UAJDn2
BDeUQgMUrcZdJjRHMKZLJ62AUP40ji8hzGHNMerFEbaJBTcQAVM1myBjfKnBIj3UDwdBlEDiRcOj
gB1v9tYNzWnrGVFRfE5qm50DRJ/AbhbnCVPSGJ6yP2LI8CyK2Uh/LuqY8prYV5EyQAnPE6tgs7nu
9mSJGk0etwRfmWx5Es+xs5CQxMUd4LWMo54k4ALd7oO0s647jwID5lJz8L+8Xpsed80tDDES/Htm
p7FQFLaVSfcCIVahplwhR4El43VRypsph7qH0tz7gpbdvMkLUaDQiS+5t85Ri2FQoQpLw3zFIE29
HbuivWVlG1v8RmV8RSf35QwOVwwkisun6hpyma0ECOkyNXp9abOpqhQcwAMMKCYVKq1uP6nm59RZ
HMFbCtr8ZB88CbzUJGNucQGHMxjci4qj6toHMle2OidDt7qLoFk9Inch/yHRmhh8NfzT5y8W1cgh
CtirbDqDI5waiov9jwvamYv6fgNwhI6hyVCnzzv9r+9rFCvoDlVeImnWs5U56VrPrMy4kRrYYE58
4UQOBy5S1RRoi/3SLIzd+yIjt2npIRqeye6CkQCCjgSnYqABxRR9oeJKmKqmT0fYOsXkLvxXIy/g
AHk+qfJI3mdqqodE4QfDxgy8Y/T9lsvPIPBs0lCh7I0AmVtvCBPlvWNEVfzdkpI4mtm1lzP3NdDW
7Tmu8HWHJR0ZuHzaZTp/9sPci6m9P6mK/08VHVcJQh4+Vut7ntRcrJOhNHkV2kwKMKQAbBzWLS95
mBFXFT/848849IjsuRoWbtKW95Q3I/wAfoh0+cWcadCvA+NQRBxzZcyOA9Fo+i/ObxB0DSLoOO58
dKng3/Hbgn1ythr9jPs52dEOOCOtVWp4T+a4ECRyV3ExQIdCY0y/u/WpNHSv9ulIt8/dg5ppYaf+
S1kBLK4cUpbdhPI30USNbGnCp6iNypjwX+fAWsqN9A9LvGo/EvWMPd3H5yCAVQQ9QRLUF2iRCKT8
fOBBSJulvq0tueFy+L1fv9drxMURsV7SH+OQYfSZe9c8dJF1RFkRvoOSdThwwkGVOcau+NUBkxV/
1Dc1Ehgv6JtVCem3zMfWOFHvlADD2uwgiFz7IdIfas/iiJTaiyDJGgQjdQ07OOSD48NienUvVVut
yhhgxfVZJIt/Irsf3QVJnw4cqlix75/mlxyJo4mw51sw12rQkqa6Q78xsYvmRZrHziasELFwUPZh
2fx3XE2BUfED9mW7ZpOWDvRvduMrydusfv4AojLxC+4807nkR9NqayHI5UTRcBpBjwvX9oodBAHP
8+ppZK++47Y20ZHMeJtni/HinxsfdQ2w+AriBoeeATXfPQi2oJlHcqUy6bs3hgxqibH0OcAqF1pz
waZT/9rQ6r4pP5GpEi3s8MTNptEj0SE9A42LtG2vlFg6fhItFkScIkrBGhyVA0rw0C8QBrNkp0rR
slKA0xT5wWxdqwmOz4LDJxPF2yIxt2pL2pys8DDPjklvntIbzclsEzM7LJ/0wpc9xjb9x5zlvcuq
5tl7wOkzLxKEIkYl0x/Z8hfZOaFUfzJbnkFT3iR5p1dUic0BY6yY7qLPgRDHVZGdjKj6SNtkWYhx
2Q7o62rDpXdNRpKsvCsiZ9jkbU9QyKaelS88hlQi+n3pL0opRqk+vrxpWNGse0TV7teD1yULTpYk
T/WDWc0fvfIT9iXSD2zGbQOXpy0BScKaIjMMeGBRcvw9cKUlTR47fNHEpC39+oZ69EUMGqtAZzFI
ExJ4G/fQ76M31qmjqnldmjc0646pGNsABisoK3KLHxVTCEEIBnZZ3Yv46PfBbw8qy2blfy8rG9am
1Zi0jSnA57cwZOMT+qT6DaYeNNuJOPFQ2bqzV/K6Ug+uvgrVy7kDfzxony7G/T0qt8Zn2V4GwUGl
sqK5vbNLMLOgQjXg/lg4yiPGrgLgXuubcFXdiqHKqwMQPaWadh3/hNKFc0a59H1oBvwH8eH7ApWz
1WXheu6U66Jmo/vnFPYKk/WYWVonuWB9uRTeP+GsYX8y+vxpssu5+l+NN0URYfgUpRY8S1OT40PY
FsUFci30EIJ5Ek/6j2HdJiY065W11OJWsu1kLIH5pEjk3kOZXiiTkHPo+Lq1f95q/XTx7tWWUO7D
JK9SV8lKqy8LXCbyce+PlQ7jD3Mi49tzmEhqwjoST83yiEZnbylv94juJtfniZKZrmlcw7+87I4u
5xYBfHDyyknS6YOlF9hwVngT2hPVom5evKWRcvA9UGqaqkTkQU4+IQMC8eAHWBz3euw5QJXz4wTX
BcGczJ0fAo1bcwtMBf08+fN5SXcy8npQoyQUDg21fvc7wjXUl+gsxcgp1d5Fp6+q2jEIFdDiG8i7
GyopAk3b1I/7YqUBuasjD2lKs05pT5DllkDUMotVcdgXvU5vFPwPxeXrgTQRA4iX5bKHWdV8Vgyj
/1H3GqOuwoi0MdAlU/rCbt1ybPRGKMMT6wSGOrfmmf4M4aOrEqIFvMAo8bRdW9VYPpKXV9Jk3feu
WQbSa6BODNXcMsKdGChYMdKtvOuj7KifIal/4OOsYkx5YNVqxS7lopbw+wqte6KmmKh74EQZVng8
tl6EIRY9rXhOF3xMNLzRxpKr3QBTYlrdcipp1i1yCj8qBW/lICFMiVsdGrtVRmIZ3UgVckkY5yPt
tSSBOkgiteiaTk/tAI9aJfPKlt6IBzhIGCCKSofTI/OxFyq18bZ/emjdRjdNMzd0AurdZop1X6Qi
L6BatbiYKH8cCLzAe9nyn9J0byBqofH4a3oITSABHs3xkxvQJLNf4mPjF8lsYJhG1e4jnoSroZVA
h5AFt7mXDB/RGuh8vK1L8b2JHbJ18heRGPzdqOwO25nVp1vFcWtBHWRsb7pGprwjySDBgZvi2f7e
PudzOWJeIQVXJkbTclb76lmgz/50oL8mFyi6c4Nr6PGUwNix7ylEeKnpowDGpm+Xq9hI3yg9deAU
s2eGIYrDAMfFpm3KNCRBnql54mQfUUh3ZyCh1wkSlEGzyG4gJoZmWi1IILSPP7s6eSMQGhgk6AjF
JCxEiGDvBKjLX3myzgkiV+alcON+fKUvVvVHMEVC/pnCBxynDH0zKnbot1dlo6xdivREYc4mqVHQ
WDWy4O5BKRXg46lsChXRhQ71su9/cyzCyNUZzq193DAO/ic79jZELUVCgbjNI7B/C1gLk0Yi13FK
ZnijsksmMGjAdZyZ+pNZoTUsoQAJpBB2j4lmjzPCGVfmWopkvuK4K2nPbjmT29bqEtaz1R/GEAky
mQnYTVJSMTsnpVAZ1DhJPT+uKHXtAmB8B2qbx3CtWrl3tswOuHW/X/RQIjhkxyHKSgOZA88lAULP
UQaPZZNOpUUZcvSLOowZsHRECOrdplyzPCxAxndSID/I0fYGg2ku1CSS7mGHcPynxHVOO9LAkZDr
Ay52sL//Wr/cfgDQ7F0cN8hJL44xRhuH6dsopUEd0wZ6L82Y3rjYTqBeKf7BzqIDI+LMk7JHvVEX
Y2GGZ0691wuJ+khR6ELtlyWcEH+o9USbHFzaDA9sIQp1/DPTRbuU944yDa4VwyZSI9jIMZ1QhK/O
HH3KcnDqaNn8iDsnIiZFyMfZPWy282W+OFjruKjzVBRq8V2Yxlr0pXvU9c2TsMc6N7foxST76bJn
f4n3ibKF8xJadr3aejiQ3UEcRt/WFnF6s8g+PkE3MkzeHkzRRerIhNeq4V3Mh9hR25ybawakZHUw
LCMQ6yWo86KW8VeAwHcWN0l3b5tIe4jTWG4WsW4NjqlxzmnUrEkN5CwTNFhporUVlxfSuI0OWobo
E+t6Cc9XRV1w/kGllBb8atggic10HT00hxplc0ZXAwsZH0tQ2MLAR64E3Qq6kHxflK9kTi6LpIX4
xRv9KAqV/n1bLEeqobg3cRk/kvTADkAgwyaDmubkohGl/LYU/OCRHg9knx9RHQM6JTUXfVNtUmo7
FHvvG4OHhqPZdsHvGV553GyEnLMr1JcjleUivdYWaJWlzniY0WWqPT29wWGrDD8mx+8XOenVdJNh
khXDHtBVWPrNbR4vFRK7y5IP+CQnQPhGRmO+A07fme8wVcKr41TqNEnvNbB5oaOe1+Wl+msnmb1F
G7B7vY6Hal63XGoIsXmxciXi8FhWSaF6KVpSDUxlR0Z6nvNEsRfs1LB0CaYpwGUQyjGLIMVG7qEW
J35G/iW6msySlRk13RgHDZrVq4Me9qX9h55N96CVSfO9cE8FlcBjzqyM0SXG3jojLqyVtpvYQrJd
yNX6jSm88Dha1CToRzOi0PyuPuuxIflhxxXNWBrd9YAKIau5t/gq9mMuq5eqwgkROsMVuH2Abk8D
9+bMsm4sNZboibcNwNEEdr6Q62ciSkyJHxULYUBpDcK9O3UUqg5wlXrszAyNPntn0EpwUhA/d/ss
Bb/0rC54kftomA8c9Q3Aa2mUyohcqz35zwrQ/hJJlzWuwGZuSxQJlbneu1bvx3H1QSutOxhNGfeL
VYk3JbI3Miv7+EGyKiWQnj2nl+o7Q09Wp/Py8ixelqFJP0n8IDZxhwGkXVzQH8jh0hDcUS4i4GDn
mRMJy4dtlSchu0P7EL0va9cdg+Qvk/pch1LX0tA/471qWAI4YV3GpVu1vlJhzIyWKtYM7x8TkmX/
uev+0U0tOIF550pTxlj9wYpgA1mlcRWPMyoTbJrCxV8O+Lli3OTtjIc8DW4NhO0CcW+7DtxvApqF
tSQFA0rb4N+D04Ni6/y2R+87Ka4RmWgMW0jZ2fTqsB2z8mJNpcubBxUqvoNn7ed0QUOALkRDtlaC
CPo9uARm3p4YiQf5rlIaEd+qoGSb5xn+xu9zDtZHet4DlesOGtQ2crVHPNK9W2WUWTkaBfdJ0CQX
Lr02xVfEstgglMKQ9likuVa+WwMJJyOCVhGla1V5kBfxXmo7q4d6lBEHf7Mb4jBRC1AluArOKpGG
W0RVxzWO4iElbsbN1++e8D7vC1ds7Ih7TqLk+CjaH7e/iam0wDEQitAzn/Ubie7kLw4ck2BHeCSY
ZctnK42JPIigu3aw6NFPxtjJ+zhqHYg1xmcJmannygzni6OpmD5D1IWAbNKG9/WPBIa7hM7dAwwG
/UKArSXIWHE7TL8v1X/CKRJnuPbHWzjh3AeIHMtYjBU0mma2DHzEdWxoh89u/QLtBs4fTSDoMY2Y
8VS8FoG34ZSohUBO+qXkRtjl5BPnKrpaqcaQIgkcb/6sXKS2K0YdmSqJqBeQHohMLOYm7JR3NPQy
mmZ2jP3n61SVylUPn6nkJlEgPO+L/tX39QZl5yfUKhc1jWuhz+WMN2JvYoUmhp8Tky/4Cfv5U97s
KrYvGSQhOwCrn8UeyeYPUWdMSX9m1KPhLkVGRB5EkckF8uJMKKjCxxpfCvnfAET1hT7IRwRUw3vM
bpDpDhKT/WeOA2yBPLF2RwBrKFUjmz7gyB307P36tgJQ28qW8LrcCU9yPBaX5Kzw84a7ngqsLKNe
vkVoMpT3gFpN9lq9FFjEaLOO8zIfB/JX/N/CGWqmHahd1OGEDu0eAg+pZr9f/NeHjPWRUQiECsLN
Y8PGvKC2fcf1c1pRZpkt9ChDLxqdMTYJeFU/3fADsoQtMWhB+iykijFtTk3QhHyV/sDoiciqL2o3
Y0TaOiLKeUx2c2F2X8607GNpJMpNAjebVgL3pjhLZBwRYJvv9giCPIwol5OrfbiMn/Y9RUbPqHvh
kFFSb0rJg91Tcu89mNJn3lOgOMo9Mh9kOFLRaYjiJ9fthgjT7gMbRTYhZa37yhHJPwoLeSJQgkYp
j4GxvtyESEU7iVg3r9OGoeZcZVMau6KiEdntHDer8loPb9s1Ia1FQii2UacLxP+AdrxuY4/Wbhji
kQJJ3gEjsuM+uq0CBP/pP/quMxCEZpddV/IxcLTITSXpf0tAklVuR9ENGS2JR1q5fYXnM5vR9vbo
95iXRnf+JSe3KBFXOCyNRGZSWL4v/EPLW7h5aSQAs4PydBxZtDKaFWNdH2SKfCN5JS4IO3CIPgPH
j8J6pqwO8A/nUbrBDj0Z9pwUMMvA9Q8l/5EOLYPX1/cSO6PLSaUqcBUXhNV5QATro/n7dCgEGgle
WHx72YRqIGpJ+jKvn31Lu4/v4Eh01tEDPRQKwwZFj3CXa5i9ZPMXwxJ4qE3sIaKgIlZo/Ib1DYCh
c/ibfIHwYTi/zY26qXLGbj0+dpWhM/IKUzsjDFIqakL3/MclQV6GKtqUoFsOCIlX+lCwwBLCNO2w
Sng1KQjLjOL6Aa12dYv5/LLsTx1UxuMn5G1nTab5g8OvNRriHCYk/7NOwyzplkddrTJNT1saOBwW
GFWby5bhSAC7CGywRJEqg2XoPb/K8RjI0pUnqN5hjhw6G1l70BjuXEkI+zcNIBFuMO9OqKvw0jDG
zL+5t3r67H5Biv70o9OBT0xyOuoiJNEJFX7tS+597VwiQNlURtjGDIflufvG7CwLgAgJRbesur2p
wi2O//9JWP8BVnz3wPB+cPtSAY88xJdCYWJqcVtEaYbSz9U0xG0HeEwcK18jJHHDEF9/45YeH99x
6IPoDpNF010pmG559x2QirJGWwKMAUE2aYjQSFk2PiETxF8iumP1f94MWx3VpgXF4HVTVDAbUir+
pKR5RG45/4O70CD6eLLq26zjFiZOJf//CR7l4ecJk9jo83EgwlOhB5RfFt14N06Zhuol8ShvR+On
eZMDbgzHj36wTpiyLyItSTitDqsRgH+paELLaiajS+mz1hRoSMSbB90qqeEw5EXUcb/1Or0wQKyl
A5deQZx/RObW34SUKS8ZNlJoPQn4KKR+1ruPpGBVUWgvOKOS8SHti7ujW+1uG4jNFWs/trmnhanD
GanLt6YqUq2mpdyiRdrdVg0a7hzwkpG5fodlTSXA1Gvk6lzqKPN3YXMbhmhbpNDhjCEzORy+XYr1
rTRCAB386DyhmN1PBfgFlnXHxZWv7mLhsop18LLxYttlMDW4ZV2mDzlBc/X6AL/sUiPBnMO9y+S+
inY55FWSDmW7wDVS5CkcAojxvtX/I8dvXypiF0n/9arhzsWDTH4ZatOfbRHygUzQEUflqgMk2A9Z
b1LDYYcNDoqFGCWRrO6T0VdPVNcSSVhdvVZNlpLhcCgkK+xarZjk42gRojgiDmbdwom/0scsiNXp
Tu9gPuhP6VZkM9avam8GPt0BpQ9Lv/e4PG1jxUlIHfuyQ3ArsMbI50goKdTPJ8/eLvzogggGgHmT
5aBCagL+A9ZBbo6jEykAQ+vyYVkX64De3YAGcrLHEbWFWg501XdDfota5Jt7Tk10M2p4rXGh08cZ
trYNBpbip9vBW582CDtpYPiiD2jU45dOOp3qhRq5RRY1vH6jMuKUhgDzyX0Zpk9CJlNLhcYxJsen
tnSl10sZ3dsFwIg0hEfMvdLYjGHLdODLmZ+Z7AKEfMQwxmeToSag8VTL6zscSCPtEnc+HDtB782X
u4jC5qVHgRCIVat3/8SYk1ALXrEqAYgYXj/aNnKz0Oz5wuUe0t1EqNK2urknBYJUuVAKhPWOYcKI
yM11sU3giCDAX88ovmrOx7enLHDzfzR6booqh9JCuH7Q2hzVBDx9pgmTjLhbIKaAsHIF8XR9/Qr4
pWuxrXbXA6U18zqhDofJxPCXO2Ra7tE1Bo+FEHm+987rkuxtQbwaYe4d38L4YHkDAaz6YehFvn9z
oqk6hq41z9mSpdogasga3l+7+1Vws6DYY7SJ+sQYkG7V/4CfevLSDTVSJ8CgCX9MAZteB0EAvz2P
WPcAm94lwa9GAfuDUz5Up+rrzsjj4Sylz434eLwb8dG70zCvdGuHJmugsnf1rfQWLjMT2+Vq3GVq
JRSm8xKx+CG/7EZRyAdAR6nzcU9/+0kw4yI63Jk0AQveqshW61yFapKtH2CSas6FvTDx1zBMSCe+
xSN0squBwEqrsROH73ZEoo5tVxOOPluKomOtmE9KiY/QWfAhI7fkGArPNLYdx2Jq4Xi2fFuHE8db
z9qlucF+xPFHoNLWdtNGgfNU4kKIWeEGfbrEyCP18Ka4zKRZ6kOcwaWkqHnlTlqmqQlwmmxOL/Ia
ozGAzG1LdCluTHMXaYj7fVQPcZdkSfXgYHxCPvTjsW1fH52Omy6SW02NjPWuAEnraV1nijIrJEDd
zIP0lxhMg+itSXOJY8VOuUKAN9YzEguahh/Cv58iB4C+zP0up7XgJVR8jmGml5FgLodWI4QofAV/
ywfH0ZmWsWoNgGS4ppq7bNb442MzLCVIkvPUu+GfjzVoca1mmDjsc57N8BQXjUyspGm0oh4E/vXt
aWtnI7LjB5crnzNx//pgNRiF3lwN22M3JzmNkwc5rQ1boTBI4HrT5whq54VvJhYAdfUPuXRxHski
FKuF12KZeVrOqkm2tvwy79flRFwaU20eR75qtwuyyyDGAC8kGf14eifhvHzlR5sO0RpCrrp1i55C
9fq7s2HBVPjz262ZWfT9B2zO6VNbizI73cNHwVaZERBbnU+idPs/I/DQ+bDJgMk/NyWpUZi4Fgx/
5eisPubnzx2e610+Ovl+4vjR5tFRmXEYnJBNEd7/0hcD6MAEILpW/ybZvA7hUJG9hlGrzo0U0jbw
vmhwa/9fSKvtCX48+WzzqT4lYCZfyHUvQj8FxIBFyNmZiJYz9oSTJgaafH12xTba4/FfgO1g9Gu5
U93WKhdx+5PODn985gUfiTAfgfQsw0Uo20Yeen5j5AfrNR5z01acnbh99EeJltFzXHxAQgGqKOCw
rRWIetSxEgQJn+Wk7z3typuvxlzbGx7ZrxGaRI8eZr0zWW0zZSzFumxN1z9vuhYMl68J3atd6YzQ
ytLloOE27FbUw/3RLWSOiPUQ03m1DwXs57kKDyLMlhtEGK0WiRUl64v7YxwjjyEJqNNzCd7GVNHI
/QMMTXpIDdGqbU+Fi/YW1BvkpIgKrkub+qs=
`protect end_protected
