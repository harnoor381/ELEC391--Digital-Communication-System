-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
aEiYDEnL62tXwT1JsRiFrYgamBtJ+zsA1Myo/7kmCX6NHCwpNNMFqD+Pr5xf3i7RVumNTlSj2YZ1
NGg2fw33U2EM8jIYXbx5jbaayPrxsh+CThsX9iF8haOnm1UKTQX6v84A3TqHJeSs47Tjg2PeCWsc
ntLeMlhUBX+G8r3B8YYdRl3TxwKnF8FJtt0oTAPlqd7B3IFyWXz1qFJMfiJEuuZfAvucKHYlNlV/
Xact20nCT7pzvXu1C7brSrn4cI6pV61Ovo+JeqNZEWr67bRHE62g37CvREbaXlb6GNI+9St08iB4
L0TTzS3e5Ojb6fdv28JJxDyIL13pZe8dGDSGBg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 75680)
`protect data_block
9eREPpgwDpWAKOTMv7lJY2FwNX3eyr8uUgynI86Ojb0JzSW4vdlDmqikQMo1J6TPZUe/nzriP0ib
KSWIkRuiOBkYHT9hbemCOulh7/1mJ0TfWPBXWi0tOsKUzecmhdDbm1HmJ7K7j02Fy4LZAIdmZM9Q
TEHiFKMZ3vdAi4m7by370NBJ05GGsNHqjPbQEURqUD5S2Myu2uNhD96jCh1BsSzEa6Ky1BeCniGJ
/g9VKGVH8+3o/42qpbB/PoiEgN2nVeIe7Qvs8ue1X+2fqKZwJSjXPc82JExiwhH1jz6r5Iw4BsLL
jhM+8OgJiqBjk/B2dO/SkhA7PF4gu2lKMQUTcLQX4OTAet0QhG39R5niDAx5V4NZKDfk1veUxcwI
Sq+FkBq3zNEW4ACntaY18hNBqE9rBlFlqUbOZMbxW7EykytKQJoOvKFBa7gkEHBcKRmRmhGMrDl1
JOZLy9dY0xk0ejX3gSqaqwRhh4UYSC2kPHPCuAKfMjQzuXyIdK+dzn/96RPkYnk+onU0KVbHIjRt
WxUsgKFVEjST1CIUvnAw3d2/C9u+9zGX0GvWDyxYPrvLEFy+7rJDcJM33YRiSvgRRQ4qgHosgfJx
xcKHZNZJyIZkyUmA5rxRS9s2Id6pOobVm74yTeYcTH9XBdVO/LeDdpP5mC3bgUKxaZA2P2khACC/
jOR7o6gRSjY2lvgSkBT1pvPEUTATzTeEqn7F2RKxF8zhpQUWl4Git/03CI+OqY2g4znlkyfvO/1L
h6M2GJD7GW61bKJGj9hKdFJXls0KR2smqcGXrDf/aYRWAqwC/V6fCqzSYgCsSq6W6MIIfPrnRk/z
mJA4RErPW33tcXOjiuDNDeYiXQgr8bBI5Qz8lGuZLCIAN/W4kRCjo6ztIw4GcjDmE0tYqVD2UyTI
MC44MNQK101zi1OKwhMEOPspYw5wqegHMpdM5INziYXXYokbyiQreQBd/bFcHF5Iaha/IgK62k1W
FRYcredCk2X8FdHDem8WjYljLjtwVzVtNaCE7+cveU7KWDEnJDfKKHg0MJK31RpPeKYCfJfw2JHK
OlrysKh71w2Zv5afexmKgdER+qKPcZlxqWRWzrFXhdqtg28h2tdKvZRdbP9CidENUUkuxV/2HrH+
fcWLYxXGX4pOrvCEZUnUrua4WH+s7Urm5ul/J9z46c71Rf12jPp0lZjlkJCNXbstEAFMYNfwxZf0
dJ1rroGW1knbbpU+d/1khcxRqvRR5uy4oa345HMrQCUR9/t0VhKtD+p/5NM1ibg0B5JDdRFLZ3ul
ChLsTEhxEff8S08OvmvXqgYfr5G4BHZFCVM8eVC5odkkg0VL1MNMaMC4Ta2He2WM0wM34QUB2Mgh
OPSa7IWB/KE8qYsCCnGpBIyVxb7/r4cjrXke/9bdMIAc/ee6e3wcHbUnq58mzlRpKdfgZmo4tXQH
muNt/zGoZTFxyu5IJWTQdMvAQnwr42w2qowvxqIxiUuzSKvhj1Djiy+gMGPow+C0C+DiOtv39tI8
kLTw44LPktBMrWqEywXtgl96lTM5POOz08OX1VwmQSCf5LQR/k1bpC5/hwhZj7yFSYwnDb6VCGS7
xQn6BFPEcF/qHifXrdC7q4Byo9hiJdfGzT00A4+TOAKIKgoMOYYDQDzGr+oUcZxpXRrurlMeaxz8
fdRFiatsAyq2G5haSaRvTSwK3YNnVh5ppmdzcswg0UyeVpu6MqMJzYVCOxB1ufpe4lkUVfYeU/Vd
rPnsrsL3fGug+EqQXvwr6UfiPPSXPk9SBmcezw/3Vb2mxMHupKfPc8QF76O7lndS/CGIk/Us1+QE
027rrWxgeVTNQ8ogw5AIypWw/NQpBs6K6ZlcZFQtsK5mDwek+k44XUVxTKB4J2dY0znLsuN7RZh+
uFwrFOZHrprCBPogwDGHrFIqQpHyFNvvSbQtQX2ZCvIskP9hE+oeOfCzQ0Zw/MV2BvIPjcLhsPKm
gVbbHciVblC0kB0RcHDKxT5zOCuOEAO0OHcStdJEgcjhHtUR9oP1RTGbajNXappesBUKcomyj2ZQ
INu9ZcYYLXdK0WPrnUfrHh7j6tSEZKQIIbT9z4CrszAsumfyFcOqk1qLUEWlYKgY7RW4/8LJJJPF
lpRWGn2eyhvWHlR7vA7ditlKqM8MQ/xQJpjlwfxNb981vQ74g43aXRTaLXN9NGEb3bEz8RnH542o
rf7zsTp7jwb5kvvBs6n0dr/As0y+xsd1OEkD9LEqn+h2v+bBxURXXpYSGEwdRS+Gdd2SgN0wId6a
19cp5Gf1qn8lKFhjr/AQbPma4M4z8Sh+fE9dwdzqJgetd6K5S7FtD6DqOFoBILngU7jUaNlYzxGY
DAZFQpiP43nXlMPz89kCUhB2Oo8s+B7tKOQl04X/+qKZVjVtsfw+ZpcBKk29edFkJBMOCylaBR+V
HWCh3T22RTvOqAoGVe49vR48wfLhBMoLs6yngGUfgkE1KtZyRUGn5/GWgxWC2+NPlIXPatZrFaLL
ixNL1m2SS4Y+WJPXuKNqDkStoG28v8HLlDOzAYAEgcxi4jjyHFgvzIsKSQtThdwH3SCk+cTLDKBu
KSIqLjVz4l5wzNH22y8ax77uxbyJkq0pEZp8b769a8EpueK/GuIeqNNJz5qQT+ez1uViVOlIN6vA
wu5BXNfSikQqyWt07vW4E6+8RqD3KBsoR8+lEDgDLHNKFkCcDUhhkNsbBildP/JDJREovdTHkR5j
OXt+Yc2XbtHAFP3zSUlogSY8vzaFSqiBd2AXCVycR/OPKQ8x7drHtwsXIryb3tBkA4tIXwNUSwsZ
sD0PdaP2yFp84/CFCmAlXbFZ6XzfQ6HgPLlfUr0mtkkIHbBULvTiRbBwCxXtxSnMeDrk8vmQ+d8j
dZrWLgEUngg5RhhSWR/NU9F/hdAAep2HyJBrHSpNeuxGxrK0k+BV0oh0fBvPzCl4hERyDX0hH12L
timRsB7LxAhvcV9wSm0Dj+ZXB1pFAqvpcxh+fErUJC3D0Tnq6WdeOvUFUSN5Nbv39w1kfJxGVaXW
LeC0feGL85cennGLbSr8U2zWBQLZT6mCs/wRE16gny4iuk1DgypUgkHSjRtslJlIsrrPefjvgjb7
07ZfhETTQ2UDcaBHHC5GwEz6N6HqBFrdHnMaH/jiyEv2970xWp43Y3K9ah+PjKiZRPUGQzPVjWi9
0wwbwnVYiR5awUGx4ChBKMhWr7ij08dhs0g2nF4+rz7nUsr+8I8JrF8AniCcZ0yVpG6tcxHD6NBs
IToWYIsiCsaOoeh55HpQ479mpC1HL2Yw9+tlQfdWmyagQs07mEXocM+b8sdu+GTgXpegKxj8Wuzb
ZbZ6TzzCnSv6JcDawra5iTUyyFb4AkA/TpFDsmZO3APDiO5keDgucSji2+Ztg7DJTOEgYIYQFlHJ
4yGq9BOdt38iRRNQbzGT6nf3N6nqC6HisvlSQ7kuxs7K0RSXAEW7XVD8PBi19OX5kYeXg0wz8S8E
MRlQbJ1D6zyxC47rPm3aeLeMTAaSH4/MJtA8Avv/e9w6vpAcPeCfSzJ0plY6moTC273ukX2WsieF
NsZnhChjCb/AS+5bnIugH3ufEx29jeQmQFs5qwZsE2ortG4i20pP2UKEYL5EsSSivyFe7hbKUkiJ
V+kAWcp/iYcDBY5rmLee2hx3/l0hXQ4+7t2Wuq83qswu9PKaErwrTzRreKj8VBmay0fdJEieghFO
jz4YBKWHIHE6CQX6/jEfh+Qb/DpeHlsX/o8Qmo2eM+tqAemICYDBmXxoPKPO5ACARtKvC8Bna/eG
3ISiHORFcErl62MuLVWE9Wdpk+n1mnC60G7/8rPAFH/YOkqCJZTceROnNgT0A1OWbApFQOSAG1P+
v6DP1X5pn7eYtLjlmW9dYQ3bF12hE0G0YT5MMMYFCAxjbxoxy7jsfQv8T8+wZBW7zl5tdhgIkHiC
63gb7xgt1bAziumoTtdWnT8KXBEZK+CMAv+o4hzojK0ciqYp7HkiR8jcVMc5716DXTMnkj12I8hA
UbTDUIHqWbNqwSP1wBVSo2+Q8H1HDvX9dpPgYvVqnlUvK2dSleIafGSa4NteEUrL+58+qLCp3XwS
k8ycfARIzJaAVY8UyzGfwPaS1suGacRG3XEoJXbCFesE1/bdpjzbm9/qYPGa9YuTxuNISgiXVEke
eK5LDnI2reu2mxyOFN6l8Xo2WQpjZZrYRP0jRHkomSR/3oI9HKcYe6cduyWdoXgLczha5szoHeMh
0nBIkui0bTfIV8KU5VOrQTJPGwc4aO2XIrTChoVLjyzaqpYJuG1NgriuxU1fhIF3RPYPNZtZmRO/
6OBP4RHdHpbwx3gRTzETMeNXwlOPzg/Dr90x320Ya/dnCigTG/YkS5k9P9krVuutyXcJj5TSGxdQ
7c4Z7+7GJL4iXZSuRei8Z0KW1VBb6PM2aMoeihfAhsnkf/aqTvvGGeaE9x6GswTrOZXoK8Nyx5zR
qBZQyAk0Ji7AubOh5lab10mE/PNyW2ULNJ3KwHtFyfUWU2KGkPZeXY8Lo8ZilG2GZsLOfOj7XPTq
nZ74uHhVLZezCshCltqhxRLbd5o+tbvT4GoSs4K3tIgZaFWJHE4tejmIGWSoM+tqqTvXHX/4Mvze
eIWtduS2adZvygBLs7n0OtTpMktcdJu72gJcG7rWUzf6skwl9jUSgnGZxYHN4niCXJO+8EcMz/Tx
z+z/YEcMHLFfLUuJ3Hg247W8Fr6qO3gaUf9+UWlNvr5VH7zcfDzlPNsI5gVnN9E0SWlq5bUuQXfC
9n0RIDJ58pBCx5hyKyWFP3aDhKgO/mkjTwORu2YvlOD47YsRV2Ea0dXBvI/sEr6xCdWchHKefPku
Hy4W/uoyBg7LOHfpOWoGiGOz9CsLkrs9Sa3NHmYOW39RI8B/kY+9nKJpMr/4q7Ekye+D+0yMtrdD
2cTMSO+yNJyvKKD+MVzepLVOfEF4+SmIGjgILQkEovbd2v5Fqd17xFxmBMfwDCT5Wll5XkKtC2aV
OU2drMTKo8cni6NzeaGYp0DDYjVbZExg0qpCT0fiAnbx3jFe1AzGI6bm2UFWXYQGa81Z9Yvzcq03
Nd2x4wjYt57dXMTEWfLuKInrXd1u7voZdcP/KLCQ2vLWjopSlumrp5tk0D+URaIx7lx5ByUskTxv
z9yqKAaOVmI4/w5sNMFTtM6eE8i6s3WeoHRWru43K3ovPZAdrk8GEWNq3mba4FlAaMLALZNZHEn1
dd+sNYHiKhWX71TeSfw521bJZ/CuHrDKIlHnJl4W7MY3zIS3ITmLrX5UgbYpJu60rFmfL7lmV9FE
AIii7lPEZZ5WgzKLErrqZscbTjsfWCdDRbFS9HAXT3NxQCPnnHjnPcZCjBXjKrP3TOvKC9tk61nf
2oMV+5Sj0opMHg6IVBspAs7Zbeej3P+1lr9EzxZ+lxfxX8SPfhAHV9vWDjSN5dM7HQztKjYWUbAB
+zF6CDvyOsVrmgNj0M/w1UGN1qdZra++m21Y7QS2R4TlSNiuBVlfNGQgndyDp2jDhiC5Cx+yfnI5
FmAaRBlVbBN/Krs9yWusR81LsAxzA7/ClMBO93jhQaOgNcETIxYyg2eUU8swe4QDLzDFQhZdF1Kg
PvzIFHhQd/m1Q130y7WS/8ucegmj8VtGfRF31K/c55TISfVCpakifLUe3VAg5fNjgaNbnmDH7zS2
g4HDcNK3mJXNcjQ9jeDpc0Pki4TSESC3XgbadaBJ3JNBdsr2AOz+x8ttXbPR/NTReaOeuHf1KAOA
Bkko1mnvVEThRsLREjLJzqQ4DATzhyw5q7J+MIDgAYL8RXaVGf6vShnVoDp4IMmHP3NgXeaVsLB3
MJELMOHIGymw6XIlKkr2Yn7p4kRcaMl278H48ykXq+xGxsYwSTdn12VgGlRGH8zSqHDr4OSwrr9Q
ONee2ssh3zFSqk6Y+xrojD6yahCl+b2N6Y2PR6A6yPKLiJKWcBxH0acbG6dN2y0o4c/8eUcZ71cJ
Nn5AkaMjfhkxL0B2qzXOfffGlJsKXTko0LxwRRmrIHh1SzJGG3QWD3vixOtl7lNKpodvxcRjQaU0
4QCQNZ3n5PpL2cicvc2zXTMdY+78NU9OmRiEl/PGmyJsbodGZ90NcO3GgEpYwHxYPPjLQD/GG6Wm
/GvW9NRsS/EJ0QDNhCUB5DuOaFl3zsuncPh8/rpbJ0H0rUyU6j5cixSpAMcAIN3i0BQI7ZT8OY9H
KmeXl3QwfXI1yf1wcXcD2rx6OH6fG+bfzSHQqfoAm4Q9YslBVJazrwrIKmNBUsqEOc5IU+QeNoyD
GpAc/yNoid0yvXCA5gndSr+bMQ3KXhtRAmnLm5fIv4Yr4tdFAVWk460n84QZcjf8GmaYSMYA7K6H
3wcEdQbbwe8AhBuxP+We6HDxI6ikJOoNqNV0LJOEq+R8X8FO3L+0CIzlTVXh8fMub10XPkKDvzNn
qWt+E253XbYABTbn3bpYqV7jb9X0xOy0E/i52YPt5GOSYsy9g5GCrBq6VuiBXcHI2MJEaNP7+2jU
R1NEn2y21lAAGFgGLt18zK88c+C9E59+jqj/v225u07LgcWc4czN7Djdge7pNQsO6mBTp1jvDu3w
k9CAjLuh7EBBfeUJmBK5SkVtTpRVkeKtLesUBLBXDOu1juFD11gdCG3+PLHYTM8HWzYrUa3jlbo2
eEIkKTco70pxC/53Tg3plI9IzXDLI+g0zn/+VT1bMRvLQkwpLTZFZI8sF08uunWAI8AikATortR/
n6HVGgyX8MZVZdLXLa3GIG9n6IaSs7wb7sv0NauEkwsh3b2Td/a8idOcTsN7IV3C9fguLa8B1Wgs
UFaECozReDNfeOLzWnbyH1CeaXB4058IUj391mdR5xcjg83aOqcvATNTPnP2LFi6KXGBibQjiPv7
+NpgGy4XnfYZdivXKy8dKsBcckmZ6nC0enRvTC5dx/ck1u9QFGMj7WKCzb39whxXBm6l7I+cqUCw
EaQ9hZ5PO5vbmQGzf/ic9sXPGx4wlOEvYqtPrmyCxfYmqC/6cRvVxYXB/vPwcAwPw00ub5H+BJKD
iu7DweVM40cL2v420FOajEIyBirFWKr8bdRktp+eoSlqeByvVPgfiRJTNC4H5lN+8gxS5+VEGjLz
oh4gsEhIXaRNqVi/gjdrwlnlatN1DjRU2W22yMklvdrQB/s1h8iUjHl78c2ygOU6DQ0BCmys3NdZ
lfOpwEJPXrHALdsoU7nTHTSWuHnkcEqyG3jatackLD1yRkDaanWfXtvcyiiPfNKMcx3R3no2RqRH
IupbNpodDYb2Drc+JUl1gULshlXlH0v/h+M1PaKl4Na1g8sgy/WCkmXGZnpRoHl587zAszQ0phOz
4MTl9p9K3l4wsEQ+ma55/rrWtxDoT3KDlirmyK8Ng5uhm5vi7B72Ol8Smbqrzx497Ad6oQozXjCP
myzrD0p5efCg36FPVNMVdNzXHR2H2qYQsFCdP4jU4oPqfNbCjPaIxuOnjeWt+7/GgpEQqsp+3cZu
9m73k3Km5q/UV2XKwbKj9cDbTBT1+Hv60Rki8IGTQIKOJulAS8BgRYyXSPElumkhH9le9KJAgZb8
EezyM6Qj4oNPKydEh2jHX0WJQhawYvDsPeoQvjyNWLKMeFM2QKz2BwyUEy4uakZv6rRNcDtcdGJl
8wfko2EvSJPugIHuglW6DjMOLrGe0vF/oLwX4ALJzDPk88npe20yb5/jlaBSlvboFgjL7vtIXwRe
kLqpFmBgsCD2NNd2yizWFpHt26ClAyg8VIfooaKhHhJV3q3Q3m10QK8Qf8pNbdlwbt/qDPmABdS7
DgRzQ7sYLPmdoTdELUDaV9eLwrLsArBn08Hg2yvJ/qHcNuHeSkX5KTiZfdNKafwLmJ85m8L5mCCo
uIfAS7kf1eYSCgZDQ2QBKPRHY0Mz+CbHW7MNmgAFkrBYuhxhbmEiLmRaVjSHrqOngugcf+Oj6HE1
rRq+BjvcfJHJCwQqsI+/ibuCPMn3ZnZWh5yXUTUHVBlrTspTARLK4SjwlLXPzciZhBGW3uHC24Dm
1/ulMMvLXQXT7Ev4wj5QqBRF3a2zT5cZP00p+IbPUz5HPBXAQwd2t+z4DMeUUtgig8wW+ZWqPnCE
Mn/bMfd9e8V+riaaE2Z0Q9bBvNzm8W7nblHiGl4WjXAAWANKPvfUZ88Tuv0FHVzaFGYBk5bo0h7d
Dt2XlrwqL3PAKGEo0Tv4FPK15dJD8d/of8T+llECYo+wODXkxc5url+EYObJ2BjuMsjIHlpUJEB8
cq45mbAiGCf5aXmgB3yTA9lUvYvfvuAeFfxIB8DOmDj22DBLql38O2c8sfmW0FU7BMPK3ITYjC6q
GMG2eaacb3G7ExZmxrNzAkks8eb+wklGsPTxe/gSKoQsw62rbDkirziLTkYD4UuumxoeoHFHAgsx
OeJqtplCuWl2E3b6QRM+0msHtl8j/TV08U7AcFFxcOIZGK89jk4xvm/yxZE7UBntzllsliY5+5Xh
4cDBV0PriUizw4sJi3aVLbxaru2wB1T5R4DhYRK+TGcooRmpkW5E9sQ+jui+P6BFcaPY2Y8frLeb
fsjkELl2JwjCIAx3hq2gFH99cA5h8pqEKFYbRurvMYcMQYe+5AuFcALaRVL6FAAQ1j8T0w06bszf
iJrVIDQbd0xIgajENRPTu6EEQ8EfC/iDefOEnhHulXZUV4nnTRdp2T3T6awkmZeHQJ4jjPAhZDS1
2sDLPMVJfrBdyEeJCNsLoJSfP4JjhWOleEKh4oWwoJ58LenPQWapM7cqhWp+WDrTztE7W7HMmm5t
8Bno/Ke55eMqSsoTMDgiR+3t6LDSucfnadVIH7SkFO2a2lSqcX1nWCizyAYlnF+MPshYoZsTQs46
SGsF9EFbDHazowjetL8vEQvOh8cqOH/jNlSmuFToW1lpf/QIfaIj5bc1loTULpO4jFVwhd+LI/do
FbhalLJ4+yuzgfNXVqIsW7FfbO39br71F7qYnS7CPhGZDGCyG8dRzdvBTFfY7Kzbz3sX7/3XJPBn
ztUr7hP8199ZLUjXnhsysUWKDKTkzuKVTIJvoqRPKc4T+8Ggxk0KLAgF8LA6hNbs+8TE2nCIEoKJ
igxR3lqr9RjNfeWd9nhY+oVvz/BaP7jHsCb886lYaaKZUjqvMfAKAZ7Ax2GOgpjiwyJybja4JjYy
sb5/cseyB/fPn2igQ6lklt4x7Rg5SU1hnvTrilDYQoDpF6MwFyCB4leQa5IVLBSYDGcSUcxV4ZyP
no5EKWhEn6D8N+YlJn699kDI8DSoSl4AgzuIFfJ8D+cbGgkK2XWZaIIowektpTveaOUBtgifVj0J
eXHTH/+iK8OkcLs89w8nltEa40+zIaxkLOXrOkm7Ul9dXJA6C5L5RdziMmUOvwqkEx1ZmD+4CnMO
KpUZRUXZBrJey3lXO0b6O95MZ7US/evasUV1pAKkuMzQTEoWp7qc1JmZITExbQZg2kyiJqGKl8kA
fC69NPd23Ro3fv6vmcc7HL9ePV0/6uzlLyH2aBfOl6gxKceBn/5vXbX/4jGoS8YOmEh6PwGWVwK8
7v9ET3nhqTWiEc+ZnbhlW0Vca2e3insnCEtxSUzICC+iwEBGj96JBtTLgi+U1ZSO31lJs6ZWOmmL
ZFgL94sf7SDmGloAkbFmQ6XRFrR+sSGsLl/VNbDWWT8tH81W5i29U9knsRvxzJYI5EuHAVjltOjb
j9Ov6zk4a2rzC0sByAkj8Km30aORT/ZuDebeeUWm9C+B6BNyofnq6wGRE9aT+M557XBLgriqBNrj
NuMLZkOcf/Z+KQtGeecz0+AOwKXNaI8k8naTfn9NxSGI6jXngbK7ltSdrQGVGOTAYdr/5jSwvY7M
MfwA5pYAxTECQW8D7lt/suSYWfSzZZB0uJOWAyEHPn8hoavb0r1gLzAcpLP+JkrESU/TZ0CaqsDQ
1PPbFXh4xfAqgSBizRXoantJsW3GLTFve0STWty4hghF4FNzMVjHfT/4+u/2Q0h/qpuubRJA5pBO
gN1Xo2SGvE9OUDs7/ZEc12c+/gk2qMZ4we/XDkeNES9MkzQIXfoAZ0wgqHsrh2MD+u7ekTAH4liz
vjFIv9Vq2nZS8VEOxWfLHKauJHoUzuEq0lSiD418ofp42frW19YoiPVnwGVs2cpChPxa+32+9vWX
rbhVzlOKpnba25f/YlafYEGhUd8/v8e/nZ670EuAs7zgvhrQXZiKdIP6Xqu1nYkfAemUV+GHqAP3
2a7WFWas37iYkAW0xQSLqGCLRfY5iUuwQMOOR1hlN7gyld9DHMTgNQ9ZaXPgzYX//0v5Iahpg4qr
6iUNlWMKZqAVzV+CYI5x1LsZVMlwMpPaq+HbNNJio7KnnQaBgg2YDb25x8h5yloKRWT14eIX59Ev
DBERCNL1MmkW7KNk9fz0k/YNZ2+GRoZSofIRWOUFlUz/sjec3l/kOlCX4Hc3Z5nDUEKdDcUH8ANw
tIEx1F19bbhl+chnNjMTeYVfeoULvbggwM5juA1v1bG8idh0RR3mFea+sJKgr+koeex2nNeG02ug
EasDEAbEPcytLFoSpdeOxhVBE09cjYdiUYirq92x+1ocyIUH5sRclfHnaISyAXymCmDOo2IG18ku
fxIP5J9xvqhUSRaOplWWyo7ybeaWxcp/WySOpqOD9YPWyY2sG6oHMdyurEEBLFWZT/n8HS5CvB19
hE8ua9bsyutjVfzzi1BBP4IYb9Vx0kbHzNULMAbiXH6UNdIfrTMvP5/9kI7ZIv4/mV3zPOxEm5LP
EFiVuRTqZ59BfWfoTmxwU51LDe4oR/KgiHkmfWATVO0U/rW7LGB9UxhCZk8M5g6UlwZ5k/EssF11
37R+P5fD/QuYX8nYFatKRnbqkQVO+AN/HqtBvtK7Ak6JgH8XYiHPtaqpGICzm/BJpuYw4QreQygt
1tkb9kMsXrZYiU1awzioxTxe8LDeLkOMnRcHkXfYiFXrkwFfFJW8PjC/LU5ZvYHWb7juYdA7PbRN
7drOrU801adpEQwMq0v87JfLVB1kgjMMaHRuIlzn8JSkooaY1LbYvDQwOFbMWC4fWhRumn1kXE/K
3U5wuCxFzxc4Crg9JrUnoKw22RPHbV24bvV1WNVJaMcIFXFEB59Qo0HkmYIm+4W6T0lHgQGEPIRP
1CyrCl8VQniE4//a3+OKTprFlTt34x96mCjyziPG0cezOcluUqlTC00rYqnIQ/ObvwMU/H1AgICa
xioaRpImtk4NY5AyKcGfrURq9zalJKoFKOKlj+0CejdBlAfCUfPsYy/0FDl8oDW+BxEsfnwHpdpq
83qdpw2xKM+0Hh8QnHhgd3BsTrA56AtaCGhik7b78IzYIctklYmtMbQatGMIJjVrMvYfANJPHCUg
FAd6bxCfaEywFc0tcs8hYxWqFXkwI7oFfPjoPX+JWVDHnOmAvs9ln6FGTYKhMlZ/42g44+rpBmVK
5H1kYUdKHL0uRVO6Y/5aXSY77O8mPr2olxnzfWaxalEsVNVVgTMJyPfkRO56fxCIOOx9opfrkw4m
0dmyH5hHkHtmfpJuau1RVPVYdaIQFHJWpHPDoadWLeC6tkV2XbHR1ptYUvYeciUlvYBr0nPn6PKj
TFtrxyNwJrWHNyKNHodn8Z+96nk+ydF/frjFOZmHeY3eemLohsDgdGj9sbRoq970CLUH18VdfMFw
d72rHZSbu+xMWmPOABHopQnPWQqUQCMLUdXLdhR8xpK3Y8HhV2g8V1AfAPEBmsPxshzkD8bQk/R3
XeCQ9uUGtf9/hTZQtY8buZnKfo6a4wF36eZHeAUOe3V9UfN5OQUjcjGoVzqsQluy23qclZb4cs/B
DwJ55VKiwk9GqRcYmHD1UOJPCYwbV4v1pb8vg+Sufu/U49ZB6caN5nhLY0p5z49QsVlfw9YV11D0
j6HxDU9XRZf71SK+Ung7FA448rhK+lxLm+kWnijrgO96FGpvKTukLw43r8+1Zfg7zmEAMsVSG4NE
tFdn8a+muTvd86/z8pL/soVZAGzpWcltNfzovGcFFJLAHNYdA6wI1eyPwt/H5oq3xpuU+7UHsZ4i
GrmqUxswWtwhDTaSuBXvZ1388VubSZ9W7Ss/jNYf5D0EqzX1sAztTIEKSh2+lQlS9VtC4RbAjE+o
qaIrEF4CJTR9FQRMlMSp887gO4cfzzKs9HGZYaQN1BzgXIZFxTcGCHBrnCeKkoZgZ+O4kH3mpExP
EcWaI1mf3gSohcMPKp65VB980Ph5IbI2GQaceW3yIDCO+t2m4WM48Ju6YS+vtSmved6Ls+UUpfVB
rH79O4U7wG/XgSW7XIKyhOKo7pNTCPxdoNV9E60wGjI19dCQB+XaMqil0CVwd4FI0IfY68yLaqPl
fQA34J0RJu0sk4oa1vy5MAUOSphp2KeAhsWtRgl7Eeupf5sWSll5CoAFrpaz00Yhiw9g8FCJDOUy
GOcfKbVrfIrcxv9yVU5YrWMI5/AoLoZwlHZguL/kfykm8aKgzpgnaD7HIzbgXObkHbu1cA2IRhQm
Vm3RJHzcD8k9KNayGXVeIVwdFUQ2mzA19PUdQrAGl4CCIp2i54lYl/xxhwGr81MVSHrEzT4CXTaM
u+vhHCjxHICLUgk5/m4FeIIyu9T+G3JNoYhJSxVpE4ehZAjGnRKDiow0HgFGX30BDvXN9qfK/b2h
PwpWt5j3jrJ32QrBA6Zmf0GMtvmoey6QFeRk4hGMW/LDDS+WYpzyfr8Q6jyanRmC3uTatfgnhz/P
2+/ftJJxJxOb8eU2rOnmOJsuGJOcDBg1ehuqM7C2qNumWX18IGIr1oMpuLaML5/eXNkVbaf3NjvX
/xChsxMPnxl+1W2OansbqgBR1EzevfM7aGzec3Zb1mC3vkKkBx1x3KpjBJUstI8KvDb2zNRPdYPU
lonv+dR+CxQGzuqxBR5QYlcS1xYDTE2Q+6C+P5a2arZcETTf5E7huxi+iw5cvbsFzlvZEs2/wr53
gSeZsRE5rv/jMMEA+fnxiNf5T+v5aNKc/JnOAuCAkjeH6Um+LyY1rW2B8IhrrTF+typORYAM9MeS
KfGqSwkbjPBXpLfQP3q9GJcal5G29rS63BHzIxrnYCaumXjRjw152GehNaIOQt6/jp32MpCsLr3x
mB8Kre+L+0EAEviuQxeD4pXWH7jDNinntvfQORv1q/0NvoSTHDdi7mYm3U8s+xKoAENH8aAcfwYg
/Uzk2uMOpX2W+mI+kRIlWrok3T1NKURo45vVJRMFUguasXEjKNghjaP/alQKsobkz1uM8qeorWGH
Ulocy3u3Ebou3zugd8mi3G5nG9ldDXwiOkUrbM/T/wgeW1ELScFT1ssm86JzznFiG1RBbBrDCk9J
eN+egwH+YQ/S0lJbU12sewmufvQeBLFpCqF5ZIeulSyh/TMw1c/26WbGmNbrzPtKaZZ3YDhVX/MN
DaYB/IUOMKqDKjIJ7z7Wsq5daz7+oITgwdw+7YGo+EpDAXgGZgtcnq+IkPH9MMtHCF2HDe+5s+zY
kppMbrGrBG01N4kjqrDBgHCVO2TWee6wjHnlmIkn6weZk6D3o2BadZ5bzaNC5srCwKW3OrLXDdlO
fcYRgel0X9VlIQbuWV2EuXQCWlcDS5L+DF1IQbpVO3gwp2Qap5lmSKvxmN2GuLWEpM7zHwCw5j15
M17/cvI4XNk8w3ONI+UfCRYIF/Elfq0aHOOBTDwjdmOMP5KBwIOu4oXdyqLkdRC4iyQEhlvtQNTP
/t30awZe9dg72BLCcZfR1Q9oiFAihioov3MmblCZWNQJuJQvKrNit/TcNQsjwG2HGkWDe92zKJfC
mZ9qNIT1wCvWwCVHk6kpBMQAa15WvQwhYHkaTP+UpQcYcnv2bSjXtn+bTzZFLZ80J4WWk4UdsdAE
vsSTEgWVNmkptNyx8Ol/HhahYKAs/VzZoBEZxmBMuhxsr06tEGcfi51U264CoSfom3Yjt8gOqerK
uL4CDDks4MyIrse7FICtb3STg9xrsV2OYOsVgvhxXUudyD+l+omj3YP7OEPCvpXYaoRnLPnIbEsc
mzqDOiAaBE31oso5utHdBKCGjXb5VO+zfi6tRwUnwlKURebeTuA0gwFUYhvb2LEoM3+UsS9D+/Iw
0Rwwy0lvUuAV4KBoIX+TK876HqSgdPxUQb7nA4TXeMpOo6SHdhu7Ehsd/3QJ2Mfhtm4cvvWJ5Bcn
ubh4zDdeuRoAwpVT/IIKW5a+SOrbg31fHybgwCrN7zBd43ffaFjs8OdRj1kZVOxB4gNjH0WJxVIr
FARXhsp8IuNfOyUgGufLFtt2Y7DkxPBklzhJ8hMH4vYh3+7ZEjaBsOWxdxPEnGclkNeCka+f4q5J
wP09AjTD1HjICnXdF8y/gdMdB8wSmkDEC95e1RMMZOv64xEbfZbqNikh5BPCS0HLgP05LD7AQPzt
Xp3Cd+wbEPrfLz26vOqHTQbWz/KI28Yjmjsg/8jz1s/ddKiLmJtGLeF6+7Aokwe0yYzS55GZDPus
vviHWu9gAeqSJ4ybRXu2vRX6rDSJAeAbsY3g04+uXeZOO5/WjOqN+kIglZbaAn21nbnySN2iGfb2
VYswaDSSeED0poeZ0p1QDV6tjrQnpySenebVj1sbDZj3wsQ9tAP+DfdYJ+lKFkyIeKte0verT3kM
4IAzxPAkV2AlOTDK6Eruy4j4rtiu4Ik3Wjoa206Ypss8OgFrN1qU9JpennzyK0spE6MvE6x8JSzM
0/i8Bm8zM+48HcnZD1xTfelGAgG7wSR99tF8og2SNSw+6KCNtxwyN5dQZDcZK+eOLtRrpF3xkQNj
jwmXUg4q1ClyVbZas5rcOGhs8tXD3DARJFgjTGXwsViUwfNda9sqJxJoJEyq21z5s9vZvJrp1Myx
0pNQudK2sPh3vWYGnoOAvL6vu5tnwBQB2dmpF736TJEmoFRT2GzWWMjT10Ie9Z+4J6opN5e6H+lG
PXhRTGVD3/oeFzNIqLOOY+9nZIub+THtY4m5JgT8+civK5DA9MbU1ZOy1EswdyDdKyQSVQBJq3Go
old6YWb5f9y1HixJKnmqc2fFCE/nA5CzYBcl7DOBSIW90Bnqs9SikLGGI/TeQSAHknZ+aiJOU2QY
0NMTqkYMyjyquV9diPjTpmvDKF5spSNrKSJxr8pYQsF7GC3Wp3arg51lBXcHT48d6dVCyXnBQYJN
BO7Zqof/3PnaNBmQ6CewXktGCZSX0lL5J5inrqm9Xa1U/PKbS05i5AEnINVgL25WMrhdy47Yx5xv
2ohu0YRtZ9YPMxcaFggrnmcmQ++h21fpUDctAuKPv/2tXLAuap3aWlJnsgWw1JmSUQbeu3hXkEJD
dQwf7+LKqhvbVCo6ukTcnxny9hOigUXtRQdCSm+nvdeSg9DXoYH+KnaOiyhApAtFEuxfbsC3p6G4
cmODu+g3ca1fUADeU7c47NuTEbQhfbpF20eaIGdnV0WeNqo31kJnXyj9mN8FUVCgyfpWjFIoyZpm
9xv9aC1Dr9z5ctc/MBdRfJFmf+zymff4IAN5fR+5N2oDyXoAfKgFT6Sv4S+PamGR4lnkotWOPZ+1
IKi1+vV+uJhQqZ7e+qpGAw9HrtTW0lUk3GBBeRIh9Kxyspmsl3NWk6hG19SCs4vaBW3W5rEEFlSy
Zp/cNrWL3h00k1bDDUlOVsztwQiK523GySNqNOxBbHbhjNRs78DUMsQpitmTS2PSdUggNsKndZHD
S/0xNAa3/v+RVXyCz8z0rVAT51hrcSezvt1/NV+maYJWpmO5Q3tiiuTG9Tzl033rlZot7XdUDY5C
IF5j49NOkY+KoWdvIL4PP9iDPsmyu1DeXhI5LxS8JdrrgKGGN4mVjHUc0gQFGSYKaGnNxbycctTr
Hq/rqVwRgcBsZaEXH2cReOZIvVQeGWi9WNORrGUeCGi7SwrlpOaNLt55Qmhx0UWFdtP3foB+ULtX
YVVqu/W9tX/YI8Gh0OJ0kETYLnOpinqN8kNlZ4hWmIiiXoC2OBjHyq0+vKRYE6Ai3sDVb4oe7uL5
wQ0uX8bmlsQZxUxzrXKASD59JZdadGkX230SljAGquvlxAUkOygEyh4tGcHbaeiT4I/JgCY/f1Cg
5TvJKOhRqrVviZJWd7v6lps8wwe9V491hjZc3x/cYSBNh7xVkW+4ScCnp928hTWLGvrgs0FbgEif
+fAJkzJOnvG3XpL0X4gZiEByuG6BHa6NE1Q0qKlP8TwEw3Jln17nkBVnd2SWa3ahgaP/rRHNISuQ
NePppWZejfpsM1AYb7THSuzc4aMzMeGSJR+exK/q+U8j8JkDuW1ZJogokPQCXik0m8kXn5OxWoC/
ax5s1yee8U/73/FvhTYHMyY284+RSNUEXRq1b9DHBgCfcVzw9rk8vdZ5U8u+ieHvYyUcpR3A1L4q
sScox6Bzg6uf/9JBRiwfU+jOuVAQwbF8x7g1RF172xUEpcbhEDqPZ9fnF0Q833vzrV+UvIEcbyQt
mdfcwtK6eE2sLLuCVryRQsTk2FSleMKrHfnlAvs42MigSlSznNHIMibkeqRT3G8sPMyBiormW6cF
uvoDtUTB2Lu2dbycY1AtSiSKtvvQE6+CdRp7ErP3ktQE0ueMTDRyu+Eeyj1WeNndZvOq1iOUQGB8
XTkgNVtlpZ58lBZJZMvCau+onIS3AOqKkZ8b0xqnPi9Apb24pB8Euf5DiiinlPumvSyVlOZN6zsK
oH5RBksT51SEUcSUWF+0qOVu61ry9j2IvQB1jcV12x6089XQ2kc3SePHaOYcxY8cZzSckEh4bd0A
T5V6Ig8kPtRUwhaoniz/VjrnTWq+OetU5mTLvmgfbnCeJeO+3BZUAubCglX+UMHxl9O/dTSCgiEZ
VW+GxwJeFRCMGV1PMWmQvWTHRBk8P6H8TvMBUCl8x6cUbOw2hRZk6PVaLZ8m36qkg9FrEXcGHXX7
u+9BCM3S6owJEVCVRofZxoUBeMbz7mcdcoYm6YC2WqxlUL2eIk1hw6CBpML9FMHofUpMZTqIaOOW
9WO+SsGI/66atTESxt3675VBUk0GdeRhQrErKa6yGAls1F+1WkWFwhbF0XMuStErN1pTUTR4Dp3+
NhkFEZIkkVsdy+55QmLhMl+1jAp+Jh02FA3+DrErqOF009p4J7RhrS1L05wtfnRCGsPQHHmqwTvJ
oAXwpLmCjVfDzy/Op6L8dYvAjmUyL3pmcD3O8DjPyjyh3jdloYruh+rcms9UfSLpun7bn7ovLzCH
Iq4ERa1t2kjyZeVj1h9WtZcjDV8X3FXYNeUFEyzU/O9OnnRt7t3y4TEJjkk0TA7VW/SJSHbDdTbQ
WsP1ZtuWBk2bi97ghlP3stwZe3Z5YO7KdXFKfZKdd5YXCTrTIO6h7s3SLylf1L4KGSe6pOzKchvC
pRJKJaWN2v8nW+L/lUBvi9Yu7Yg/jHH4Je7eEft9CtAbzjkKbDjEXM23rnHyNISmGEBPvyQR+0VE
pGRfZYju1TtJsHjzwuZ1jR91wJg1tlXKN4L/qW13DzHvXZVdtDts0fqvVVq6Ta5z69Suz6C0+UGi
YwRLyJrtViCLJZNeepZuJlt1A1CqPiYlz2Ey5jAPxwagRxuKM27wDXWxOoGOZLYiscNG/q4LCJkk
JzyF1bFHYzB8kxlQRpMUBxe8BbRfOOh44RkK304n7Umh35fWAQgrcr4gGuIJgs//UldAH+OSpn/k
gix7VrkR+ZzuobepwPl3ObuIr6gOIzTHdm6/bL/EqjuCqLBlmSFeeWYHUHaXkKoZEIHGG93gkKJ+
jHImJIdkpsbBpkv1Q+efqYftDefprDDnHLiNzwlBGn5g+Z4sZr76KBs5XpCRinhc80VweKJxagiQ
02xPg6pZK4dRyQ99zCg3qJQY8kacOp5sLHIllw0UUpfOdBXZuyDLTv8Yr+S55A7UKW6d5pS2PuNo
58DycEL/obUUKu/nHDCBHlY9HZTdRz01qcIYtEUVAV1JvHzEBqUN5dNEQAud06eeX6y8wBaOqXl2
Fof11Of99DglBSM9STt415vDqG6SWmFFs5UlDePVw5ttY2yiczRdOjTA/gN2W2qfyCgL9xf3QSQh
8gGhE3fdmAKGqy4oVmHNuRkMHKjKpaWO0/raesRbx7lNya50EPHK0JCpXSvEBIp8Zda8zS3W8WyB
UbooTOPOu90pct54KCRlZ+yTa8gF1W9UAwjam1ojbaJc11AjjtGFimdHcmgCZpA4/XUNOJfAwupI
PhjeAReMLl5co+/uOiIiFBVMH4ippJxphQbUgwQ6dO8OVyCOdI1CWjFE0bRKQWmP/B/LYhBMSuzP
fXe9nixEVD6hsPU2OUfAAMAAH7p6mAsC5AumbM8fSfRSlaHTsh+Z7w30tQtTlOEIgY1m9cgpYpYt
Ob3c1F15w/zAmNICNeJlyinA24Tv068e3p1iMBOz1Fy9GVExrBA46SED2qNPSJ+GtkaABbPLoBM4
MsILa5FBBbe7wETCXAugbsp44Tq+1BPrWIBBtfgmnyQGqEeOwbcjPps0jueWgHw47pCMTmt5V0vT
pAPW6QMfKQWFiI0Z1gRM7KtdbQDoncKPrPAsTg3zvvAcwvUAatNE6RYk29OhoQrokFjaNqW8qjwg
+UQpbZaobjZjlu9OFIaSorORO+OFQDEvshQmYZwB3Oy0JrSkvAjh+T9p+EmHOScYpFigu+hvu3Td
a8ii9Kk8fu9BoREbvGmdV4jLN9fudtn68qOID1U2ewSrFZzYhIUlPvI0OwnxD+0Kc0UWi6pSDv8o
wzvDXxSopnwWrDoL33t1+ClrDPWrBq0NoGOZb92Loo4YqZ7SWXKWV5UBR4Y5nhY/vlq8zznNskLc
On1xudg1rSY3MnHcdScH8g7vs+EqK2ZEBgC1b0fCIBxIO8l2kN8jxisWWmDa4JnlMhCcdHN+mW1m
cyRUg3CK3GJilqyheLm2ve78GuMeE3pxdr4ssB7IROGiHNy76o7dgyLc0m504JgtUB1fl5RiC1OT
evPB3mnwR/gvNcZAA60B7XM5dDKqUsUwEpil8/NW93uIBkzorudrFwnB5+Q8cVh3jq1k2LMiPbg+
b2tPyrBAB8160J+fpgOs6F864R+x9siOarkfD9NeLxLkCu/JN3KkURp4m3iyHFNk4o/dRw/MmClw
HdWvY0MDFhArLQwfQd1JKtIwO5FBfRfiUkbpj35Ea8nICRw+jtLcLa5TZTXcpNI5XZJHQFSJWiyE
NQkyNC3pUVWdRiD2FLr18vW9b0Ohaie3TkcX0yMwaVRyghNdJqg935SNZwcc2he0fI7duZ4MYNd9
P5kBNNSIpr5wws6hEBqBxa1yi1PKdktyQEdHrSo9ApRJs20Ogg3O3APch0C0OiFxiXqcNwBdhz19
3quBvjYxnPbSXSyP+r2mb1UViHQo034NW5JeoquUOXRvto0MJdY6ZJG5F9TavRt6tBZQdLRIqxLz
8wECM+fsPZMfMY6EZ6XshWpz6miComVYZ09UT2DJOuqQt9hsVYkqX/7CVA73kq7+D+U1q2LBCwVc
SgHeb4/EHWuZQ+38ODgxXutt5oAXilt4LYM451A0m2uAO8f4rwiJjT+PF7/QnAwDp1p0xpxZsJi1
0AZy/4cetu7K4RZBmTyVO92sJoN1mSLtnK9ntb7ETos4DE4pSJEch3nKVXMzO8UTXtRVY8Tlu4aA
W9TFyC59OJ++xm/IQ0u3pSW0+POOu+of9kGZD+Etak4Y6cKsXLNHAaSLqCt3aT5hWtj+tcgsROK6
pS64NN6vZG90t1Q4SlTM4kmbKpB1w+5dzv5JlouIWog/W8OpEcY8cNz9XsWqPFllJRVvN2r6vQ4v
YAfBWPeYfqaNGvNNNI4MYlIEIR5ufWJLCsOpbvPYLbEsS0BNetfUDCH08+dwCnUCfMDpAEvw3IAu
zvwXBTKdA1U9ZM3q2obQxgtvfQnQEXm8epep1t2foNLVcrRBJxA2oOHoTnQL3UMUX7geGy+6S0AX
KKF6kAMHVd7h28WR16LojkXITwMtOVDtRyV3Iw1P1mL8dI2H9H44nLM5wiv2n0UAvejpTFyO41jJ
iJqXF/A2FNT57C4TwwZ3whhpqZHaRRYouT+EZ59xzPZyO+Z0xqL8809Ikac9L6lImLcgCuYWWYvz
2Xp/yMVEA7dGUX5ghGAjj81iimUKng9yK9Yv15919m5a91fqVn+qxDKN/DVP18gbBd2UGuXFE1vC
QsU9K1xLZU7wqsNYgoUkyletr9n3rK429x7sn0NRCCDybBHXI+CxZ61rAiC0kg7RfIQnKcG+ozc8
z6dVd3kBy6dbfhQcFORroIyGHBzLaXZvbX+h1QEBf00ySasuJpj60o+DU0JDx+V+LnmkMk3kDnfW
BtN56IX/NGekZx/zEm7Mf7XnCIeqdtGBum+tNskFAYAuZ/h0N4PqLTYm0SueAgeq70hUhbhp/KcT
GHO3ZP9S9mDZmQ617b5tgqxmBuDC/8xIWEPdK1Qz7RsoZ/1F+Xcz1IXX08zGMUkgKqdF3YRh7ceu
oL9gC1PLOpcMVWJM3ZXetREisUU02Q8yFMsu1dheOqgeIw/XU8dWG/oAXwI1pLIrGdgDRWAg9uyF
TfPlVXcGy7wJiywU+TcNqkun5cteyePQN3nFfx+vbA9hDEYCxxZlcT9WkUusUF7ptEQQGl4Q86TH
AiniK7jFZpIz7AzXvRq05k3gBHZLavT+K52NkAVhMkIa/U24OS1xQljkJnl6WQmqDxb7/Rx2w37f
3abliJ4SitTYKws9b4AQUXKbQ0Ubu1JIf2Up2LreiqYiCBtmJ97J7mDQN8NvhGqLaDZbMRa1C1G6
r7k9RfNMR0rDaA8k7vu1lKm9r2lCEJuRzNlCmFyucYTPt9ZGBsGTfJi05ofEmYqZ6JqOAVMvU4n3
FZzXmhgFdc12yXxbeUXH/QE9OL5j3DK8Wji6JHjV4drjFhDTLVC7OfbmQVNhCm0jgkDLYQuduiZg
FrCvVX+zYYl1SB+rsLH6ByKNYWodZiHmkANJezaCj+1jRPbmUZ6zYj65SxwRl6mxCaFyEQ8ygyfw
AYl02VdeX5q2hs0p2aIy+DSurea3Qk0Znpdl22hwx6e2GfotCJyzJ0170bAsanfAKsOyVG6nLLLc
oz2/hddA7FKWry6Kyi1VoXbGeYXyjPsFKUDpJsSfdZ7M6f6Ma24mqCAEaO4CHy0wJh78QPBu2kUb
4VP4Py6/MWR1rHgi+yqxJSeNbBLzI6zX0KWzsagEBqUANgOmsjjamE04t8o04AQDOgx+wR17hfEc
l+pde03l/Lpa9vwJ6y+J+vRapfQOedPsJ6fr45GuPBBCVn/8qw9kAA6VYyzOiQNjL8M9rU2nInO3
rqAdjj7FOj0c4gieYWsyUGCNHrnBsOWuBgAl2gOndJKU92vVYpqrPs5rU74Yazy1XfSNSNRW1KXV
2IsSayUgecV4RILWGzbvGRGZBaLxYCfRp9CxCAc5SikiDsQVaO8qduLl0tv+O8M792kte3PHF738
A1MymiK64eOvFlITQ3K2nYRaAasTNK0+UQTa/hvbTR2eRt3tbEsgHp0J43/VpAx2Ell6ugu+p2Kb
fnpJ+xXPxvo1+E/JJmmhHxwDLI0LOD6GFUAYO91inAKRhkX/wkqMUPpeTzLhkVEQVMvHE0MInKoR
cQ73gpQuRHr8v9Q7sxuOSxGySWJcSwDR5TRpcoba8Z4kpqfesF+GsjipEFLUtR9E0YJzFoHKiebH
AJtuyIlZrpAo2OFPumEPFqsYvvAHjhY5jem0dUzN4YxIpQeQ3jYLrwap/fsrVCFl3tOXXVgtqPWN
2SpfNToHp3uifQ4LE4d7uo7KG5DaW4/LkoOJNr96WhyVEFCWhtOf6f5CbofCPZJCXu7YQmS+eeJz
5a5RnWt/JwTQuY28hJfWcKmM5d4aR7rtgTcKtTIFrctgQx5w7p3BG6M0tMa2CAoZok56hR7Sc2z7
e0lmbMO1G/DmLH5dlwJDvJ1m5VmPvpLQ/KL9ZYWRofS4LT7JmrLDVeTn7WS4xYWpSZ6+57VUwIxk
nULtyTIXxpcYr+E8i7oRHSO/3XNbdmB4ggXdhvywBoE4c0plbTDN0ivTz+RgvZy5I9KdNcfwnUv2
+cqx4lC7D/to5UFAht80RHRxj7DvDOXMTVGDvpQEh2U3Pc2f9GA5Gh1FOWgpesaEJl6OIXwQsqks
QTw17bBdNYO2ZFobAXW8mQUfLymm6D3Ilq+wc9CCAkLgJc0Pn8pdIae64c7GNzmz+V0HmztdL46W
FGXHr3CNMJ7hMsA8jpW0nnmXf4YiSG96BzRXYScXZsfR2v/Iz52wuQVH7BKrxJPwXcI9tMgPi1jD
hSkxgQhHHByLQTOPDZoUTcfZitLL+GuIZfP3b8p5cgSHtAKSrP+xUGifYSkv3nLxZkC6+sS+CZPX
E+PBdr/avrVqC/hQpwZj6mroTAT9ALr4LF39fonnYP5e1e0qK7hW5P09pYjJ1RSySQAnmP4doF2e
TG3todZyC/Nx1MMKFScRS4JVnP0VK/ci4qxVok9S+RXxPTp9UaUhxrf66aX7lC8gVfzWuFprzUs9
/pCISA4oT6rZDDB2sZDZDrWO8sA/RqzD3syLjv3yIUbdlqQQvEfPinWsiEREzqiBgahiCma9wgB6
hvx8h8GtbNRIEmRT6sFdVo0JKPejTO3TDZqx7cOMZu6wIFbdPodiuKhYFQexP/tGHfYDgX/m/r7U
AbCuda1i6rFfW1von4mhGc3H5jBuIRL8zkK15pWKDzEM48L3SbBz6jbrmBZsJIkkMXbILsH34CHi
smDQJqCyeW1y4PTOJMBQWTZ5uS9pCwxKw2gOFGiHY9fZpSASOXn14h2A0wAOPX8Ps8HhsckTR/gT
6ZZSxNgqS20Oe/8fmRifi3M8q4IPKhUr4Rw/aqKkf68sqsim3/1hzDTEiGIjNdSXfFCDCv8sX3SW
1yudePW3AKeaEvTjUMdYTMHXRLFAoAPPmXp3EAsvGAN0oNLojfEwyFDe/doLBX8l8cbeirStkMio
NZbR8JFF76o0+R9HKkL/CU+++UD/P5A2EUNYiKMbN4AJtnL8X2t6l7e1+Qn2vsN5z0O29psyNdzK
aNlEvAp7uLkrjVsPUoseuUYsNeqe9i8d19Xq+d/+LYliJzp0FgEwAlVPTuzV6QATr5dhczJupNMK
Ww6jLBfw5heBked+zDuPKY11Hk5kZHh7JqcHnvJKe/+PAPIz9SjikC2emBWIOHAdfmpGek/egFWw
Amybp82eV3Vsl9c8k5/ukAx8XspxG687O8b9lYVxU/LclrjnimbXRcrQQJjxSE6HiqYBCYRxqUYk
p6Tdy+jiH8P8rYtY6I4uanaNdIRbPTgmSFNLSnQlxDKU++9X38QeKYGnP8DLaJL0Y/rDqu2qN97y
9iH4ZHHQm+JwiSuaWJrwWxJyVfpakfFO3Hpcpg62h6wsVtRKA9rSLaRWWSpplcm4z2kfz+C1qT2a
L6EJYzFQC/8qnnPn/LISQ2xFKq5eult+16Qj0I1PKmfrMxIeP3L4unwjjO2QfhY0QO2mgRVebP2j
7x3s0QMRV/Chq9Tdiu0g+fFw3F0CatHz2x8RVr6RH7LSRhFh9TuFMSvh1//PiEWKs35XH+S4m68S
JHloOWehnY++1twFZTjo2YSWgLw/CQ8GWqOn4IRKmaReN6VxWktxjY/LOGBsMsapH6ToaCHCrpWf
R4VTSOvCRGZMdMrvhiXo0/cMhCKLE4nz92Fymvpz5BGkhmzblVkfv9n8Gb0j1VintTs8EJIXeLr9
Rs4JgPj7yKss+M3FzhlCxtvcrYhV+kgONjBYnB26V3YtWdhZYiinRWKFBQe0cmFXYdOgj9mePTmY
pbu9ePQkoJo1XUrvhG566mviQNLrotUBdkx6UUIbZIaHI4qyucE67f8zgI4cQWaLfwnQSJNWLUue
G9gwRyfhvRvW/vrJocYusCxiedPjWfGlvleTUd3zyLYLisBaS6ztif3+xSoP11myHdc2mMwfqx3C
AOqAzYS/t5oqEnSz6A/Ex5HCjxlt82A5jw6nO3N/fPr0RZaMecxja1pB2jn+ZnsZgz5JZmPMoGsR
ScpJFkL2JP6M/V2Y7Xow/c4/CQI74t4qUIsF9z0yVkUrGL3zHATahgRiHh5CuC3Gp44NNTPp4vbW
18KKz7Y0Mgp4TNvZMqr3ctqmcbSuTMPVuCko+WUeHEkteez+zAHHZr76hS65EgQNgqXqvoxWoC3O
GCVT/D1TSugMPrJe8hy6orFiZ2Nu6jzDuPH1bsXmIqCLj2Whq7M5Uy2/kOhaPoIao7vm6rc9p/t1
tPsomy2mGWEGThgu8EJsL6M+R3c7n+F0Eh+q0GtifaIQOuE+gdOZMAOSUwVuTKejZOhum5BCDvZD
cyij0jxDtsyw5PQyxs3Y2KLLxSfn4bBKylZ/Rfx34DaXmQCWf9ZUO7nlsmGCW4/mSBh/ylOeCp4G
qmBe0TokkW7yQE/VmXnsWzZdrWyu6CEGlV2YFuRD3gZP2tvCGHGTwX+kZmM8mOcvFHkJ+FnOtiMt
q2QLnbCdUwTP2S7Enbc3nGiwsZnLxE1zsxS8tsFtv6S1WimXfVic8CVjSK5ocNyYbLvHoeX7ZZTs
9+X/DaoU2fVq39mAXSkiODOdIxdlNGRiMMSnrqQfXJCChV3ssRRkXk7QWWYHsngVWwHyBbLOFcfn
SNuoIngbMwxrGBaUQWs/r62SGZtunav6wk8CUrE1vGrKArMPon/5WqnDHgiNm2ObwKvk+SUx/4nz
kFcThj+VR0DXj1tDJU0nrxdweCe+ZX26x2SAVLHy3Fctxq3fIVdOSWIGfQ8f1J9f+7pBpI9nZLAu
meXLibIhIRCN4wEkRrULOwbsuF10R44lBTew95f64antjcXRScR8Vyu4O0xRJxQZogyPwmjr1ktI
IkmWY+pAjFYHN8mgOeHCDd4IVBMAKcDlzJyhKy7GYWGgr8XXjsEo0B8LOVOaf9FI413mxSMEqqin
RtjKYQAhJbsRKkqn1qyVK2Iufpdk4zM5JiqZglzGm4cLc4G2c7vBkvRTuarSNizPD5uMbMh1bF5p
BNX6jfMrOcCaK4LnilFjdME1RlyRCIRI4t1h5saWnniKnX5iV3hwZWhNoryF3jH27xda4e34yq+D
FpxmSaR6/rkRD21cDEYE3dVMaSATNiiVa1vQ0bA6MVXRpUVouOPwvqc4giIiuih9USxPbCfdwpSz
QOR3zPoxEm33nKhtK9CeOHe0fsjuv2+SBcuITzf1g6VApV38IU5bQOiAW3e6C8BiGCvn2tIkpVvZ
eCG8TxNsOZysA+Y+By5Us3mKjuGjwTEke003vbI8axXO05oKWeEy0np66YjzlBkFKfbxfCZb9zTt
a7lZjyV5G6EUNhF4PElKoQh8IIlfOt9YpMKzGZj85A5dnqIDlbW539irfj7WywOiJDgKOgM7uOS3
8RnzcYDj6HaDMYHxXOJ826vwvnePuDZXtyaRLglKkBorvdL9JwBlYWSBv1tfjZj0H/gaODEh9L6E
3PaLbCvUvjPho5N3asUTuTyfcwXrV521dZmUPMLjslNaTJlcbvqSecpLuPb8CRpDOu4J1p5Kvu/+
V0qR9EtVBMo0GGq7VuNlE3N1fUnCClDikQB8v6GFk1u3QZEN6lAjFHLB01Rw7dwK6FsPioKuHuVF
0VgIl/aJXUo3bjs96hayoG8CdSIR1YqmNKmAhOju+atOMSbSbpmJsz3PwRVA7jz9nxtPXYisD2m4
EhBNdW06GArp3LZLl7BiBYxb1KKcyZ2yffJCd1vL/zdr5GGjBeQELhpstFof1IXnta2nTpaRS6O4
Mo+mJIPkzLnZiNsJU4136LxWs2o3fge+f9WAnDlN0fqfI2++mHoAVwRfOg3um/i0L6fzMyuMCqvH
dGyKBjlNSrIIez1Lperfpwv1oYFmlTeW5iLHm70QU+gHE+Y3AgswmNYZO4uMrUzm4hHsi3EIiexL
XMd+Fnv50mY/ve+f56CvVTkFViQvd73tpi/I6VN2QHYrFW5dlLCATXRa8IToIo4wWjxBPaBR7W3v
tpjqw9mUb8x4A5ZnpVZNtsJXMNoRdVKVpWuBIUN4o6g2cejKDqZX+H2kFAI998Ct3cNsI5bJ3bf7
vuWUO6/8e1dZ9lZHJev9YQ5FOeF8XFPXMSSsXbTDLE/vwRTNnLASSDMo//HgZjVV8WbDJW9MYFcf
SWrFt83kovnOukhHh9ekkBFVh0V9OxeppydFJMpr2+5ZmoGwJp66280H/8YREBQShmmIp5CjphPT
jiU1epKrgivGD65rhlcb34fUnIFwymrHugmxU+8NWDq8bbBGTJAqd2CsmH9/5SrVmFV+nrIHypr2
8Sb1oQrJex9wJqHfBTT7Ty18BiUvfFLsuNQsewIGpGxVgH+x2S4cEIAUACvDZXQsdoMgfjMJ046x
7sW0UlQ1ldHoCEmaHEHPqs6HMnpkbXVL1LOGHm19hJo5ICWcumahGFr1ChSEu6RJ+7XcQwZu1Vln
+Eb8lLdC9QXs/8qsV3U6JWoWYsGWt5GIrJR4GJSTvw4leY/BdZeTXQdRoN3sgUn6YIuoNsr3+oZD
wFcBEAkvTYrYtlHBswMHdVk4KbgtK9R5ucNG99kXCWUzzCeTa2pbQBVNlvGuZ0VjpCfPMTEd/88Q
DVuJEWYMJIF1gqEF32CelhAOBDwoTXsAMiC/Cnmuz4cZOw2D5loRL85LshVQrmf74AQxPt+ylGob
s9MTd/93AsvYYbP8sIea5ZIkjcdIsg2SA6piyBCbBkfmlZdW5YAZLH6EaPTLtgUqv8VJFw7y89ur
MWKnkfvhh1NHCsbod3zjb2Y2W7EPVf8w6M2Kyh8WADcIbLW7DnERHLg4xacHUNlvNnEJhrHGCDHn
9UEIKxLmNJEKClU0UTAenfOlIMLOjGxsGheouPDfwhb1IiM8sscciwcK1cEuQaDpFnR//PbmLsjp
ZDdnh9/fVYT4i1k9d3AmN1flEiqobi/6nn3N1wg8BZqosfG0c7Vz+4vTZ9X6FHJVPe3jTtnbn5o7
47LGyztuNJzfd7se3wTYylXEfewLS5NM4GSY9G7hVeDOOsTZOzo5zhesNnNs36CG6q+azThzCcXd
3KM26zRul/rpRhNKFsYSgaJwjIZohJmAJn1nQncCSyGPjQ7teZj6mLZQcag/2G2TYHf0ZNewjyAZ
SOm0vB8CTR5xeEVN2erPq5TAMtNmhzID56sOgNIl58hHZ/8lJef5H8kJQim3aheh/JZpKGYLvOgw
p/Q+CTl0XIOqdQOoukxCW4+1m06My720gI8qa3MZSod8Kq1JpR+XDNRgqrc9pgA3/IDZbmn8n0ez
5hyjtcQ6wb+GVfGocjg04gHS0ywLGmdNlzLjRfNYBvSn6wT5Gdguju9JaIevf3ZwAJhxzls+41yX
E3sKytp2sUM8b4IbBbMbKySXnNRsUIa3uALZepOe9zu3KmwclMy6ppejeN9rGjl8BJKd6qAiO68M
2ZEuNc+UqymH3mDiblYi4GAyusQK2+Q5Chq8EkIi4U8jqZijVtwqhWWNKNnQKRCKtXEYSMvSpuXQ
nnb2ku/qpR6XqJe7ladATCMf5x9tYe2OwoUOP16m5W3aainiftIywv36eIU50n4HQHTqI91OypNO
5pZS5aQOXXwPpRSv1F4MTR1i6Lf8yviUHcRIK6DTjxvf4sPTC4yXmRfiQ0fr2AAsKChiAhxuQfoc
dDVGzMeCMOC5sSQ9kcel6G8m8bXtqmB+XJRkdrqwvtDbd3a9tXq5L+azG2S5UfjlpUkzEd6YD1XV
B/HXV8SbDV+LdOI3h6EmqqWjuA0IAchBaSW7IJbXg4Adyvv0LfFkZHwUe7PjTFTwza9xq8c6rfIp
GAJE0bNwNrtmk2UQ33to3Q344+aQorF+dXCUA06iuI7hIw5N11A903PrO2e3PNANCpQTXAaQ+9rn
iV4jcuQoTETW1PqDr7V48jQhx1ruVMhPyPHPxJvBwVaeSE2lYMx4DEngsf5Bd0HNI0coGcwGTYqq
DC8uJKNRYir39wqXS9v+I5BEcCknrX2BNBkfVeDmjaLwABDjbE7azZts1kfv1O7wHSOiJh7LhDVT
oY7R4L+xZkBvdntR9kaJtKxfW3fAR0yrkUGa8AL1hIX+9OBv5cI5zq8fLj3doMuQ3xA+j/HXy/5s
5MztdR9eKzHv3TPfI9D8vGcg7oGCFeG401orYs5BY4epahohq3e29hIvizwUWUBZ5iHUXqNk48VT
WolIL5jM6cQ9SwuuYIaQIJ/hQIXEmbzR9bWasvCAlsWpXo3Q1UxSvEotfAFO2RKtneKrz1XMp9G+
8WFT1jNnfj6NwBfPRhB8XkZqxkxBsvy9KKZAjNwvQSuDiM3xX32U6LneL/2XbhbeMyOYY25G8535
BiCu6wVQNtI7QIxI1mnbNyFBVLN5zafef19qsnD3bQI3TN1jtly0V8L8TvcmoPDKZpffOLnu3p4p
u29+7eZ7qsH+RRttyEptL6+o3QJ9SphyOHpwmzwC2zMiI916t7ByyzX71pJsdaHjRZ+zBgYuTIaf
bzBQdcOroJyHjOIp1dqAGkuBX9FbSvvnMpBjsfPlbDwcYcn5KeUp7CBbyA2bu1BuS+dWDrWf9g90
cjm4AdWRj/CUfMUq9/1NlJjflv8uxQyrnEDPr9osOBs1Ks70nW8o0WyaL9dcVvq+muXmR14AEPGA
fkJfIZPq6lNb94RZsKUMxtIW9wz0ir4GYYzWgvwehaEPBhCkE8AQhO5VvjH0GPs9O/vDeBdzQ+TA
rO3UZji6Sd18Wio+++uLrrtR+W/+lJ6//eJ391H9JHqpSGnKI53eqGJw2ZeVMUaL+Lw94xiRtDag
9CBhUz7xfzB64h/9+GPZHP9hdnH6pmZJyz38CptfYe23qhg292gTYH5+eq+mvYDucV5UvWBXTufV
29dCLlYsQbsK3swbvhGc8QezYEpdpsWKwOV5xM8yQFX2HH/YbZDX7X/hIH/zzYR/xayQh5SUVPXC
FsclJns7ujLB+Bxk/yr7ELns63/r31LXz4kFJsd187pjfH6Y6cpBr8TWS1VtAOQK5AmksRcEqX7i
KCAtiF/sANfyXYgEdS9XnRVodbENO3JdL4fb68TRc/T4XNDigGEmnNemILSdPH8l+ekm4Z/ZCx0L
NRCyoaAjrETKPZKNAbnWlS0QVCJi9Jm3rNXdFXmlVJRdkBYZsLY9EL25VHWLonlL02K7ur+MoGVh
QgkRH0RB9Dwi+MXtFxJoigwe6EYKVYy8Aro+xFs8sNYMTtf4gkINnQsjFlFRssno5F0HtWgn2eRd
3Sn1qIZNv594iizEZtY6Z6w1DR/3hVAacREUZovCW4bXWAaa5r6hJ8Bxaq+4LvFjlJlpWbkWV/qV
hlQZirugDOLq7xQHvZ3da1t9tWSj9eGr64f0SiuB1G0/0CYsNdYqeWJA8zKfOywCODroLw2uPGOc
Xg4uVLbAcz3Kd7nEFkZvYB1WPmSK2PIGbplrHzyS2WU4ZETvojaLEjwfZA7Siu32oWc+hnqwaOXX
ly7fuJu4f/Tveo0Uw4uqYk8adJuSkcIQhTWvV2Hxx4A6fr1+xzheip6wjaxSl5nU73YO+GqEG9mT
tPxS4hVqkZ2m3gcB3glBK35VDAEkK+DRM4Ds6aHyRXl24YF0C/DfbYaZzL0LlvoDr3mWQKTJRk0E
SycZglZffpLUAABtHGaJXlbJuaH3lXJ+XO4ytH5qoJVx+hSN8rrr7ibip6cUDC7lioOxTt2/NTey
XnsEEirLVufbHXrxTT57wWv0SAHg0qOJ/3+jMCESOKwWGLAnRT+raw1A+dAbAb1ap7o9SHQBxV5n
qbIOcuuptEejmiYEawomHObXcFR0/r91A98ertxGa2T7KbhKgn2p8fn5s3DtLWsA6+dZ4LoZa8qQ
LbByuazEblZA9a1QtJei44iQbS8+MwSVAAGdqA24no+NwgCsBC01nZtdx3GRWjjZx3lojxa2hER7
GizIa3DyKhqkwfjACI+0/TCXJgCmDdBeOMhnrEfUMeYHPB+CSrG+UjwGlV6wS9Ffdcc3bT0zkgGV
W2inirVBV9wqLrlvThckL8HBFL5kixM34vOn70QlVNFP+m1jN0JwXT5lgl93e2nukJC4YmjKvfUF
u+K5bVI3F3VWiY4kYcdYoVC+0HyjZ3DObjZrYC2RJZzA+uNwzuI2iG5asDsW6z7oBTGHg7YGMRII
fsRoQt8Ysf5gdHAS5XNhidYKjOGn7xHkjmefIYiFrPTFuVAiWkVrHzZsgTfKFwvAyC1cQlkjyew+
r36R6s3+tGqlhIVBMnX+e1CxFDRPPT+kpS2UGz1LU4s4fXgKq0o3ZnMzKOIGSUviYVyQT07mE6Bj
VpkOTf4ccrxoHxFmKKiyGm2XMxJhiT8CeshQtWrpGUMCfsBva12SNKPMAPiVZVvPitE3LfxUH779
1mE3ZLjEqY57tSexD/nCNdLJNmyzlomhJeFTksRZrK4loZVr3lrpx1w8tXYzwEOPQw/p7KTf6Y39
x6wYGHfzVc6N5tjjRiBnMDaEy1IPGtCQUghOWcd8EbFsyZJ51YFnTcqOtde78b1BCuNtWLGeonDW
qU12eczmNYh3ksq5A3OTLshp+bFMUy/86GXgNtIOv4sNKs1x1O3OE48ZjZxQ4SdmXebPFGXRhYxg
Izef2wGEWqHgFNu/I+61suCj7UAURbgV7kvRB+bnQ1p1kXChCAesIsUamM0cE0Kd/tZPP0f6GzCL
E9g0dMR8Q3P1Lchv4UjjogmeTsVitoL2mCqo8ZW0MwI5B20c8iGnApwQ2g/piYQoUzEyQeLj9suR
N3/x95Dgj9lthEBQMcgo4cMv7UOSSkdNUmlUdTMRh95wkCa/taKTZRUw+pugkHfN3wJb5RP5OZje
ha41ACVqfhXsj6Is7X5je0FEJY+CVyzK5bOIGq48w/WFDGbp2vEZMcMS5w904W0VbIup05xPh6MD
Yr8H6KGuzSjur4wpjhYDiaP2MOUfzqRWGyZf/n8lRiBCyohj4nST86YMOvcQxnxOyHP/iJ9Bgrf9
Spzx6gtkx3Zm5BhgSdGgyvMsb4PKm3elyGXFg7Af1B8A1ZPMFGxshw7Ub7i2SEXtOv/pUzfriPxu
76DBaE7tMWZzNWt/4wQCmyt5WKGdTpCDezxIOirP4hRyCV1ECVZDh3A6C+pxuTH9GHqkrxW11lmu
qt1qbq9EH2yLPXQP58YizZ5lR0g61Zurzu57R0qwrhIxVEOCB5ZezJzJ2mAS5JnX7QKwyFge6U/u
8T3YmhK23kGqqAI87k6OhH+One764Bzyu7YrPUvQXbFcBctylDZNkrhCgWBS08EZtBcv5r8CxTUP
ZobnO/H+f40gwZjHhlSvEQjUM4SlyPfWZXfVwk4nNHccIqxGEbMZo7SklTIuIFkaAioBGBfQvfI7
DdKGs86WbFQkH3G/1HdHc2LTmvxCYIEk9CnVeoCtNDeVI+1PQGF0AbaCJZ+2IECUig7+gg1KbaeS
WK49uMtItrTmEP/2IGJJ+Q4JzKtpU3XTg++l244GQ+NLD2j4fidfW/GuWhrtANyWkb56FO6G/p6r
4lYAisHG2wh/+tP/OBoI105+y6bxE51muYuhrBg0/bTw2D0w7Euklj77Tas/qPJrlDsbuXKKIkHI
HdEjJDCmiiXwBZyLd4We4a36OJH787zBCzqTdYiu7q4CUp7W6yLUEkshpNTb1AEVyoDG1v92KMWI
2ONYsXTn1WTZ+oku2rUnBCp1mKpmkIPZlIJY4i4cphWNJHpiWKsGXuVJeDB/WWH9+6iyfySZTw0L
FDMbFaS7MkNgVzzYxwOVHA0uz2xr0WoPml/H+GrSS6yol73HkCMzH4KA/CqQVXcbj7Vu96LVJbxB
uPDmKTAGL5SJApgigMj2WwMAOWKMhcKccmlkf2+DDItnl0GmKcVpPjpFHrd8QTbTnEfT6m3xaMRH
5ukZsaAOxqRiD3RIqLgHbkJsxHRcH/2q7oe9xJ8OWBS5zL1uoC31UQCSsmzEWRPysfPyri/SzAKx
6DxiaEvX82cITSS4aLVMVVbtRKwzylShy4YtFAWCt5qyJeROcQZ77J3yhpnLb//yYWzx0vREtdH5
mSpA/j7WVhQLMo38mvNSJBmYJc6hFhaWQy64/YWX8T2EQcgtHY9wAl74AE3BplVlPAeLkBK/1iNt
CfwAmHomWLFE4RdTQmu3Hfj9dl9GtTaputRDtw7JaQb514G/2MqjsQLytn5P1yOIWJCTQ7lhkBfh
WHCyUx5BP0OF+1oUkjkhtM9PBAnCZYib3wD3CyZnp+O/zQfmCZs0X2MxFK7jWLxgjRG63ZkUcd8x
qgoihJz9+nUnCGjla7xu4WYwADFCh5a0sMMbtOmM9RZGCJI53gdIyE9pGhuzkz3/SBtRHxfT/7Y9
CzHYrB3kvjRPVrInzzESUhr9WtCP+EMVL4H+MHLj3/ZviFFqZPe5UoNgky+jdBMUKPVTaOeqzqPs
JIydD0S3Msm67fdN3Jz2mSdb5lZ3qanp3jrpBod/jgYZ6BpR2hgFiq3+pW/pNewz00Td3/KmpLy/
fLlnhLEg0Faujh1v9cEtaquOZh2NYKsHVaNZ/wPY06bfQ6VMFzMZOD2h6BJ/hBUeJmmOuNfUp0tt
itj4EnDPEZvQwnFbH7q870pNd56BgT1qe4KZ8TwigWNeCUn/VwanTkP643S9TKqm6hiqdUfPlvvN
r+NaR4Mn7p+aiCIZMVGFKXiEXSyb6J8Q4WW6EP2m9VAsE5zI3kPwNSn+XxDc0BZLIjPTalQLXfXv
zD45YKcfnpt/pxmipc3PF3Tq6QkLQvbQtBFMDEPpgscwXIbg7a9isInPEUAnaLBFEAC5DE4fuhL1
K8A7xEsHTjtfhmPEMboyk8WrOvnRRiUEzt0ebzt+TSkohHWW+CpdvNKtOnSseODZ7+PQ3i0G6h+D
ho64pqLneKAbMGAQM/Nwc3kVcVj1fzUBRJtsL+HMyAAVrjD9uqXMAQFt7VbVtj1J5RX3eqWnHMfG
qWl799/hMc6CecJJVr+0TrlWXGIeBHUmRtInWm9A3Qb+pxf2YY7t4jH2vEEXq3WyaG33Ifp24Kc/
SqJ4ulENlfAnbz/eFTBTHZj4YvFwl+bH9jL1hPt/b3aQRvH9upQ8tAMSkyKLIC8nyOTCecc42Yf+
58NJGFg827MLQpECbgyNsk0C/s7xxHlPFSr4/K+reCkw4MRqWCDSI8AqPqnHL+uvmxZRoYPlmrqz
p5tthPn/ldnMJxi8fEDEAmHvO4haETAFOZRVY1g2uvhtvUcR/vhsdtQN+hhpPYW0JDRyHsukJEb1
2G3Oo5VBa4Sh1qncTaJeHHn1C5lWEoSL1ZU7R317FDMXqQeK8doM8f8tsTQiwvdGtkmzpbZYDjhg
oObVcI2/hr4171vui5orVuZdRsW4pNlQ1Xd0ufDLa+WDJRwXsRPIkednPG9yEHVpR+98/1JvtvL1
aoEiezOTBqReT+V2NZqQMz+rSVG7g9Is719FatIBfSQIktw8MnzwkM9+AXLWsjEBga/kDmNsjx35
qPKC+b/kAaW7NI3d6jT66PEC1U9WyyBGjrmBqNrlmaUPVV+I+hwwivi8x6Z2RfPyAXZN8YGFjsdH
+23sEwDwWgn16AtwCpR9GI2J8UjmudvyoQeb63uo4BXonHmHAHsnqAxq0Md4PpR7VWZjWJ98uGSg
wyqPXU6Bh/DMyXCX1nqZGuUXJiFGUvBx+VW1N20oAWyaDjojXppWLmJjlDfHgNaanDghmUja0mww
g6BlC0CBOVnSwnM1QPc6K82BWEExgGmTXGPyN5Avm7StDwoogGJtoTknuCfFYKm1CgnIIQWzLg+M
hmA8V29+rZAB+laoXTqz+P1BHcSPBTePFPE9no+9JlHC+IMfjn4+LM8b7puFl7w14DXhnAfImaMg
DeorsfzzN+g74HcyHiYaNbuXD4EQPjK8d4LfIyVpQheJQuerr/WPL1vZL9hf7nRHdW6Hwx59K6OZ
CZZYyoq+ouZOsM7dTbhCbGWPwIuLMXnwtLUF+pjNSg1GY2J2sOMsoSLhcEndbDXfvSkyQ6e/7VCv
5Qr1zodhQUKKobyY7jjvATgkeVfCkLZnp3tNAhEDqe4SiH9Js88yinhpGlLbyk7aCZr6SC4xYach
RVDxDy+cc3vs+O/NQTKv0N2siCTn3KAvi6rmdRoZ6Id4h1adKsTGRIiypcUGZgchEa+2LK2QRRZA
gLtbM88pnvi/EArpZsK2QMKWzS3UrzLaf68CGuBc/47GzVE9NcM+7MgBzL+fIL1U9OhFlUUw1iOh
wQmfsx2vN1S1WqGQ1DArjjDxpsVMW8GwOc66+3AwZHJi7vNIOG91M1ElpMmPLycyZEckDZF+JyC6
ScxPxv+TnHc4IrSc5JH9QJVUTx56qPjKq/v0qz7kx1jx2oW4jdmI8IDSdooGArLa4SkBNh/ZPxBt
OA3gxVnK0rVPV+FpEPSf/lKqLmPJwDV/KkwdIUkBY7NKt+dgp+4Xk/vz6EwSkk8ub6CoBvltWuNY
Cq1iatK0iMLwzr7DRrv+2K6tSwdWFJ5hLejNswwTwGYD23nkYLryulBys8C/2j8A17QGpycHErzy
ow4qriDg2+gb96UauM/LsAwG5jLdDU1doidvhmo8wdlqjApHCNuQkOtr9WBPOKNxfjdC+fzoqWbd
ONZJAFRT/oTWf/Y6/pjXCAMUksV7w2P1ojd9dua2tVKO79z1nWHes3rKu7Ip1vY/H0rhIcuLi5SS
m9ev+aRD2qhamFP9tgqO8OziMw4rqnkb2Unj94qS8iRHtOhgS9xS/Yl27TJ7wK9KANTTQW6ShJVP
ylK2UaevvxTC7NLjmk6ZeqLAz6i+4/6QzOR/ZwBwU1APA+75MDgz7s7RnLprG+49QSkNMbHm+qH0
xVzAXEo89gfYgSCSb9r++nxuHth+K2YQGKFyJ9i3D4Jkm475t9FfQpOhZqYMb1+AuuovmlyQlfNd
OKpKCbyrOy+q6cItZhl+TmfPHIss2ENyUC/1rjemBPZ9bqpXTsfN+6RF6xhxDTXcX/7LwG6stbur
2DLm1R49F/bM/wciKIS5gkDfV62wfuOq+fnGwtOOzaI3sC25S9b9sFpYityFj87sNVbRpGflKJbC
T/Ib0JeKEspMjxP3PNKJQA4cU9dCY5VSTiTanYgUl1DioO5DoxVw8miepJtbQo5FXw9tAhkntEQ6
m34iwLuLzG7qrRoyByLbcDtjWSO0Xt1RVo0wxTb5a4MwYERzdlzqGq7NC1ErahRoPf88oMbrMr5N
lXCLC+uDxdb4ORDfLtioOrNfM21HT/QP4H3npUh42dTc5X68OPGUPQx1x7epKaQYTo49uAzaodv5
9DZlrVFTus9Zc/3tXyfYg6NNJqrTxkM2mcxZ0SU4kyvJnsB70cv7QrQowQnwfwANXjT0DvcsE+Kl
WmOJNqe3rpTD/KHgS4kafUdf1iH5BJ9b7gd8z6vNQOaqB812QIQpAo8ZSS++uZw9X7su6OUlLkdR
ZG4gZQQ2ixmwfFmL8ujsyUGERf0L8RGNLdcgg1RbOMn9dUJL0bLhnivZ04bpEV11Jm2BAxdJQLuw
ZGqeR0ADXcLstKiOAzBtDBot5TrjNgvxQQdHAq5TmczKHyFyzYw1c4wXNaMAmFc+kyl2Zr7J6Z9W
Rj5DisuhxF9t0KiX2zV9dM5A8Xh1evcxtcJc0n+Qf6OJrvlwKLnqa1DPmsnxE7sCaG/6EpCK5eYQ
MeizYZ1XMO1zE6kdGiIAFKLAmfglaucwJ6Vx5Liup3vx3KCZd+tXBhRvCMAv/n3HM7w+4ii2FZCx
VPry0tihjtBKhAqy5uipnP0ryVqm7x6I3sdob1dvVrJqLaz8+PHjdLzXMlTMWi/4Z3HpFqpKV+sc
8zNmaGPWXvpxqKCUVLEUOogCgrYvst2K6ya6BeOWA1cKWcSIpw0kzkA/68d1xKjwYTAodfbwjjNE
LW9I4uEevDfakGC7ck5LpU4x1uiB94ZvFLzfKTVs72rPZ1i+lrEm2zkU1Fz0RSwCO663/4ENeL+Q
cRcWqZXsTfa2Ecekm8/A+yWpmkudBpr7OpzkHRB5vt4nkLNm2nYtcHcBjQq24o0N1JcF48oEtvcc
xuOtI0zGiPFrOJdu4d4hlNuTcTepPH+NNWVdgSLhvERLm289NUS4BT/N12eDhiTuIU4bSXM6d7Dz
Bu7Zq28+wcqCpQ2Kfhp5V74rE2X0IiLH9IX2tsfUSgiuzVLAUyRf4xkmhUE7/lH6rSWoK1PEFnjb
8RCj1s3qG68RxHVmcqqWW9GLH0raOTBOUVdkBT4MGKVXGcNgSHhdJDQF4V4rjwZyjMuW8TudzvGM
GriTpkX0CysuCN6q6jq9q0/EmEZbTvvL9vI15ga0wIoiSQUcxZ9M7vKwPWIq13/k679flNA+AADn
Q35XNYwoI3GgIpkkmVr4z2ghoHz+/j/h8sgBeo1AEqftWhPO/l6qd0cCDWxNX8I2xe3PVLMamH+C
+YQDn+R75Wz+5q59EF8vMgcX+BfsDf4oGqifpv7MIXCgSnh51ff8IyUFYkochnN2U22JtDQhuj19
m8ciWHOhYGzaQOOo98bhFqietvN5QrK6j2MZ5CrTJsf/P8LRGliONsfDZVXVtOlEaRR3cKTMLJVi
uERt/Uu8OQWIJ+hAn+Elb4cDiB4Yfdk7FrXjhzabxgPVi+yMVScLZO8QBGEzYMVyzx6UZ4h8qS4v
/fdaGij4136pLzd2H/IG6ScdRhlH5Z7HbBtzA80FWCrvbXwxu0/b8lIzqrPwkNZBkxFX6HhxP/IR
F1EZdfLAiLWR53YvQJrgUcLX7MWPJxIvkje5rnQVjJke+MatR5auOSDvjZNanYOAE69MdaHJywRc
vRKfcDfKHsM1r6yG2p9aXn9yewQpZgEBO2gASiHmv4Lz7xWw3rtYkAskMVzHHGNet1vW3iYjMZIP
CyqAbW2S/mt3SbjPkPPbjfrQuI1RUYe1QQTYYyCGWEH2LEWanR0KjHId6XSQYXbp+xqhZGU3s0cf
waIRubx/RRYTx7oNWYEE5R/UfP11RCi0pxW9uqEn2KtDQfhjTc+JSqg8QYzbU1qZuG8d884mXOPt
5EPv+nttfq0omk/G6AlBQu6jGnbIYuJBb/LUJAnqLy7vzJMOQzzfJ8XrGzDiTmfbg3pr3fLEOHyV
v0kTB3BRWDPHgEtxZSBJUu59N56AAkQZ9lnJIIJOo77hSCjaddECf0A63x8IOtXm9jfvcVQ242V7
6CjuBGgIX0Qg9COWDPsRGLaZfOTTrJaUWsw0F7j/ILYSPMnaDbVSf6qIz3fRVpRfjWKnBBxNslPM
jXalX4vlxH/g7xQLIB7litRtUTLUHSS6m3imtus/gXolYdaywo5lkj6tyNWT9ItLrLEHNLhiT0oH
o+tSmzhGcEfe3b3KdvdN6jG7JL+kulw/fKQng14CYnE0CgaeBeewEnMN3+aSMGE1M23DbcWV5XUz
G7091q+IU0oVW+cXvfGSUrtCBcmWOQguQdVg4gQ1/Zi6I+5DsXoPf+g8KfHGZN2UhYpexS3PyWCI
xVI+WMUi3D7oRkwFPh9hxHygvOA3Su2yRdKNqxJM4VVp5Fxa1NS/s6Jie/6+Ylpc2QDjlKp0M432
KnrjWwN0RmU9Sc1dfkI0MPwkKzjUGD/NUF4xtIwxjxtbbFWqcxeNfJxbyXF0UJ9XF7gDPpC5rQkW
pJEB1ygCi0RHLvAiS3oYbrcFBX4bja7qnC/tHT46z3iZ1aMjGgj90F6Mm6sfa0BQYkZREAIyVGqF
N6Q2jw0aqe1qrf0DGcg+GyD/cZfFJtn1wjwf04qc6egNyzAL4q8Ngeg7oTpo3S4FFE2WgeKDEiXW
OcposavxVSFKx1UvKjDPpA5J1aSIWke8Yt0ruCegM0PuHB1KBf/63GsqheJfUfwsRqze5XEft/oS
42uDp9n5uSLBy5DPqy4ra1GGJwFA175QXm/FrxmonW/d6sCB9WSH5ckuy3NZWrHmlXWLpNwp8Rpt
TNNOsURbhKjGpNljZHxOFEmHmPFTXnkWZu/ZpsxdwdFAT/NhLHqZ72a7SnKZkf6jl8n5I18Sbj7i
H8PK1durTfOlBcGhdfsZWpiPmBJ1q6HosSYiyBSu3j51sS909ZxL0lN2Y/QqlsZ1KMRdmOiX95hk
WUDZUmXtnW94ZPhgs/7UjVDKmLeQ2FLqjLWjqLDMKtAKyu/Suo7wSjh70lxyM56pQzDhau80J25r
u2xh83NFaUi3T75kvrl9jkVu5G6wjTJ0/7ihhdz0odSSvhRm1L1BPSHPdMDMDKXJxOVKaPqlWd3Z
Tey0yLm8+NrHIjVgS2gUPR60EhO7Co2vXkhTIH33+QK/S4GibV/53sa5fa8ZgaZlhZ6AbuZYr7Jp
LW9p+WyoOYFE2GRoEorzNiI6913OTo/3pt3SapiK1syJYAAUMuNTjdhN2FBb9vpgItyIjaHNwFyQ
9p1vAhL13x2p/OUTJpp+cuBP6CZbLP1IqO6S0B/HTw0h44poSe5tMvL4crzhqPY3gVyBy/pNW0bS
k5g/XuaDizv/UODltYJ3LAJoIxeon0nI8ZUkmzhgFSlfPaHwUB/kfDNGUm2t2ipgEBrePtFblVGP
B/HI0Ajr3mS7oW6ngl/+t1tVEu51oUMP6PwKVndguqXlqr56oXwuNQcLvgWcGphFmXjhmhutFMqg
9cy67Q0fo+R7V/xczxACtQM2IBQ1Md/V56N8YhT/ylepYCqKXr/MRKA0bxc70jVBeyUZ7OthWZRV
7WUPpgavOOFAifzCPIN+XtrMJ+v0TI+M5393iaPKmKL2jBd65CgtL6HNXnDFqFmv04y+8CMiQdHt
ThMhk1ZCVHQjbOy9zWO176pcTWXAiQLauQMNtdvg0ctmEvlO1R0pT67HgnYW8odmXRZxdwy/AxUm
se7jyuwRYRuX1uPeGQpMyU0IegjpQ+PhCuuBis3G7wtoWUXx/7C+CMYeeqYnjpO0lhsl56KyU8BV
+dgX+czS87GnMdNoTuUzCEi/a0Cw2Wr7mxw+SwZa9HTUEtSvvRmEW07xS9U3jAhsEHV49C6P5pla
5rEmqPn00B38unYCbd9ZRmbrzxQKBe6aaSJtmUIaF+4uiBPXuqz1CuFN6vummEgYOB8bfaHpru+D
FzW3K5zQEKM/AiRDkqeDvdmRUYBofCFslfbrlDUXtuCdeJZuVN+y01GhgC6CdH+Qxf0h5Voo7KH1
WXeh0dw+yp3hSel6Jcj0Z7l+qGqkB+bzQK2b/QbGouNo/OCBwNlqpx1bmomjcDM8JhOS7cO9n73x
J1ncjel+6e+E5My13d3zNlaVBqZGIgjffrqC21Wrwc+xNnm02N2XX0aJ3GmetJmqROoqZApdGNG1
skWAd937+2C3hnWywsMj1FRrIK3/5FotRYv6J8xYZ/QGwua6EeeADPqcR5K4N6r5OFlQvW9kIwRC
MYWcR6Mf3Ti4tQv+Ms3u2esssH89NHvY8Z6DAkkdHlgK4sQBnHK7mY2DrXzRpu3Ope8+VhwJrih9
AIYiGFXAYRRUplOb9P8zaXSRq1Qx7C25QPqkaKOSvIgh45zgPNVIqHxrD2irraEa9ogTCn1yTat2
sX6yWdxVpiFqnTq2R7+Xo26NaMsCXodiU+w+17dEVbNx/EAAPtLKaZvu/6BvXlRqdRau5xg+cJVr
McUrGNVElJKqkQC+iDUhwAM2JwpnFovZyEp43NONPZdZvIoQPj0DobR54fFlUA+vz+VXQCMFUSzj
Yql88kLtTxU4s7zlvP0XBBDOFUqsa9xpM1YvZAicZD652Tl2wm9PquwiXnreXX8/BKjMO49bO2QQ
oLYQouHl0gH4nsRqBN2DQ5QM/xvAWh4ElvmTkOW+iWt+UjBFyB0tCojZkGo5MJXwRIQhW1GZbdTG
dPRiNX1QuxrEjSEhXvjPtS3wO3+iG/Q2yZydUN6pMOEFbKWwoGorzxBHJZYFmJ8+Sh/6QjWhbGIq
ukp6uYRM3zpnmwb670KJLuQNZUol2xXzcG6pdsSUwp1+CG8c11E8kUYSHIxELAdz1pBQ40+CV6Og
hylbcS+bfg0MlB4RzwoN5ZkdjRZIdHa/65Ppl6cMKWTqSFF+UUTSFPygUfstVNW/JC1zII/Ab37L
OllpFpKa/8cMlD98eyBuudtzajWf0zEpkJ02DDGAklgHkOeGoY1HIFW5JxJdU/IjUPU5W84dGrVZ
17322hgku8i4lxBhX/7/h+YDTwiCgCgmax2IgdBm91pZCAGjfT82OHBwAaaUsmczfraavo9YZojB
2rCMhLYBhKuIl+9n9seGBSumdAAG7xlAeG9nF2ZvEzPK+Ry3+I8DyV+RZdv27AAytWV6+Cut3chd
nxazhr9TLjNp+0HhBPFL8mUpc1IksYBTEDKcq/uwEOeHz/3UsSbBVAMqSJ1r33R4nS1WCUZGrWhF
KBFzEAFJswSfW+F6RFp0Qx8HEY6YIU3d+kl2EUIOZzQZ3TvwDhevDT2R1PyvlF80gq57AQwozyET
apI7pT61J6Ty/XbIZitGTgOpexG0TB+ZlQiX3mWd6WHLMnidWUvmW7a5m2p09fjNF3n1P9+BtiPt
RscokZxkbkHAW7nW8rUZ8C7o14IsyIt68P+1qJNCqMxFUvcnhsmz0gHTUHANbOXR+5ifJWB5nhM/
Z7UKJRVmbuE5ElrH+04gf9Xb6pHKV6NlFhRVIoaKe4GxqUY3GV3fByNuQGItnEemJwVb7Pn2lt7h
JpcbgiM5AmThji1bpREXh0ZJJAFNIjmE2Id0HEOkeCdKFvYWRUtaq/G5pynCTdwA+NEySsPBfcxv
142GH+6amxlws5pctilhtu6COLkRbb2Knz6FisuC+dD9w63M5UsOfhHRsnaNLs0vGyuy5+EfOPY1
2U5s7d8kI10C4oenz9bOCOJYcreyP0nvXHH3VGVq1N+NK3f54kB/JrDIUWC2IjkQebFJeU2XgRr+
Z90Ffyuvap16iFXX3u7w3NIe5WvMPHhmRD2bX1ACLcF5eTJSkBA0hwp54bpgy8Sn+jAWfE1gMyoM
uPRvgOVTx4R2tM0Ga/O03UiFiDX+0syrBM6SiysmFt0gbBtacKq3rEX/RM64G4ATw7tKv8raA6BV
se/10sZMVuyQhvXFxCgVcP+nQw8blKYhZaFc4J7YcjRf5uZyGZKenFgbFJk107XMU3ZkyLzdtA9B
kGN1MF0Czp+X0poIU4m4JZeNHKaZx4OgoIXj1GtfiHF8RfiUJefAgTbsJ9gEOXL2P2h+EtMvbc2L
fGbYuf6DTmZFyvYp2fHSklUhXpIPHxClJKI8+Qvkrs81DuFDhAbXGt+KDdqiByRtA7GwtwEySbyO
qSDZ6yS3VRnAUlcLQbb5HNk2tDQDfGrP6SP1AtS0lFjrs59nBILaevVMQwxqAUx/9ALBLNxWZbBf
w+gIZpfEoCQx9uN7IW4mIXhPPr0iPpIogsfixoNJfe4mdMo7bO6/QHxx9OV+lX2f8iuYmYycnBjE
yYd9hBOpxWiTIZYLOYksjDvnJjLOMSFdSS3ziKwqlR3FK7YRLv+LN1Ir/VinwV9PIcadCKm+ZOVB
d8LPzE03dkX4T0pandxacjiMeYuN29E2W+3uEopl5rS1/y5+p70xGYPeHd3YX+oJ3qzQsZTA92i4
z6IiEtkC+UG/XdiF1mGAHinzrA3hWi6N8K8DLsmYMV541endMfVm45uyTGZCfTTjk/m1tCL7j9BP
8rVx5f5Bb7rIJ8JqAOJYL8R5orwLeumQta12r+LtdbOWZUEJ+rBqPV93nQuLK50nL9GOUQzb/nuT
fZIJz/xDPQEzUqGjIUDJbNLeZYRMq1xsiMaOQAPgf7BJ6P0Nt9MUYKidr8xwQGyBwQ6sjAu1JQBI
s4W+xHgT0pL1qm8W4CnwiJziUp+vKJqLomDGzAI965IzmCxUT9vZVgTR64zSVoc++ySjLs0KDEMk
klAsLNqUSJ7q8ehE1oxr5ibKno/t2AgW91a1TAmhoj6E0t7IoGIx2lhTWTnBPql4QIRB9qtF87DQ
LWoactk/IqgMUeV7nTvXhVYb8Au7R6paxulb04WomhTXVvgtewFpKDZqnVW9TkehJhOU7o1JaMUv
83c6DhQTjiHDXVcjUBWFkw2IQ31OGavpqZRrlUncbP7OB6u93JLnFXG9wL+BrLc/NOUsqomQ60eM
JzOVChL1itBsmxMhndSY1mhGq4zXkVmWkKEttB3SC7DSFR16TBrOH4cbqVgy52xW4uJYWXUB6Ty9
5dSCCYhLGfRUTDiiBhqqDHgsxNCKfnDD2C+Hh11HHLPJo0A/3YHRCmFdKaduhkL21NW6ibL6okKo
ypeowbvfzbKXm4o/hiVSr/f86JJGpacYzv+f68cGBGyo/WCfJUjf7xZAC+FKwhv4sNN5ad7xvOYQ
SBVeV/1ZBwafB+ZlpQPTTrSeQvm2AydrJALuOaiBcrmZyOvFg159S9ZE/2Hr6r4sgAHjMEaJB/Kz
nWUOhhJ+Edh+q/JaVW6U725IYMfvZEYvgBXEbtRcPDOLdDbbXlPcJgq1MqcY0GiOhXlqscUEGgPx
mi2EaSHvJxPCV8ExgoAOsK8Fb88Byg1QxYamNqBaTYqRJPm2RJllHFQf/gkajrGJNXmJL5Qd+aBb
+7HNlPMACKhsT3pQcxhjnWZvXb/pm4cyTKW+Yt94A7s/l3SRutUB7DT5LYx/gJ10GcoWrNeXliFN
ZhxA+BL4e/Ks8ujvnAlsznIeBq7n6fSKxLyYsESfZqXhOi2sNSiykNRqPz3h0cmWRT3Fq65eNqah
S/fO2APv32zt3UtLm+YrSXNwS3p9FCCGHfPXwLLHfy+DA1ZHnfVaXOvLuCTv/0ZlSfKLxEudNa+6
LcfL7RxKtHaX9ZfSghiGk9uwU7Wgt7q4NVS+Vqj7tDVQQXGLWw3PVX1eWIN7dBQLhj23C1ZWaaSs
Gu/FGJ2X0ahvjSlU4BVWTGv8f10FJbxizOOP6G1ZhqQ99ZJuO1g8Yppvx1vWHrWt6A6z4jd4Tmf/
rGw4LWnHdW8AqqNlfnNm3M72VcMIqDFP9zpjbcZYIjtXbcVC5QGLEADlGmpsjBmwOiyAitq9GgP2
fkp9LGaI35v3JXzPCXHLrvFfqd2kSIx+8+FtiF0Q0/lkjhBabohplgPgnGmxCu4NzqQtC92Prc1i
jdhdVCjzgi6z8WRQ2sRNqIv3q1vUIwX1LXJK8VM1RKDIYawrXFGSw9pN+zqEl8pVTbo2iia6nH5m
U32FZerXsCDtpKsviBdUnhb8Ux0GegiuQFAAqTGzxmQnr7PLXm6CYNs64Jd/m48plkRWEyx+R/x+
g14im15TCK9SmU3z3bPsPifDpiUqD8hzBac3mQ7zlZPk4FZEmCVQCgXpUt+jD1v4crRyW4imQcY7
QsQsSnY+12QLYMzSrj9TNgXs8RLlzD4cEFi475OwTk0Z7rG+HLuqTER1558gQQa0zRhx84yQKw0o
jzgulcxap7Zbk3T1VvCgpoXITwLiJMEFrTdsd95FBIBq1FjS1RgZaJGxRj3A7UQjmDt+xf5na4aZ
kcB95xCva+RoCUXEAT3NA7bb2mFR4rwyiakcz1cH9kVtT04nF5rABPlFBjWsll7oCBfuoqOnD0nz
6DBlYQLcNW/8QTCvyFEKN2jhnoFxchHRimW+QFXRt1zmmFNPMT3Kswr4vPPqxgt4vmwyQcDR4RjQ
K1kjvabI1CWr69RUShDXfKt1bl/iZfqvHMoWgLy8QyOJAydZQtIFlKGYp5u6bPR9INth9at5Wqpz
N2cIe+83DdZj9d19AXDos0IU/loj5uT/WaTiNiMf26Yd+Y/jmVLQA1tsrcXnEwsyBb4HIK9SWKDJ
KLHf+gk8SKAAch7jeCXZxII4s35gPeB1ocbFEsXkWpOMSq40ZxFvqQoXJ5BDh+MjML8P2jmmthTi
r6+Veyh7DbBc7jXlpTWSFtVMXwV1iG4lXJ+qOPbfYbgPkHBPqL2aglpENdF80qy0e0au9Yis+Ivv
m/jAje8PJZjgqoNPSkG+4T00FlWosRBNHSkY3Wk0XuXXo4qYKLG5GlAl/5NfQry0XK4FqakNBr4C
K0ybkdI/76L4BIEF5nJk+0DqpLY6409oqcDoiF48nuFPLOvsiMi+zryRxslne438sEeJ0I28j8Un
wojS0Qa5ejr7xx/mpkkIllqpGGhDX7QYqT53MJkZe6mZxfCmEIKXHO4HmvN/junuggUmtIUuoCmv
xs9Wq7FU5AIiEp34mssjdk+cYPLLY2ZRO8pJj40URW6Xqo+bIyHq7Yf2KHomDkhTIp7k5AkKJ2/c
xWMh2OIEXMipLPQMLz2Ttm6018EOfBhc0KVpsbrzmWTg2JHLb0pWg/+hjVBAKEbc+A0Olh+26rbk
f/vbNRChlSIjtv976C57aoVpTXnqJqEq9jD8pKKlMHs+Gpp5sh41qzMJZyJGhCv22vKikhJREznZ
FDcp5yGaEEJi3DiTpJOjn7ruo9UsCHpnCmCJ7Lc14lR12NzAp89qk9J31xOpP+kFCP53mv//0O+T
bMFUzDnrZmEH1EkHXKW6FKZZK36EXoVAgcr+GnSIjOa2RNJ4RHTLIuFM4aaEFXd4PGaaB50+YkLV
BgiuvIDEOyV00Pgsf1AkVUjl6pdDA62JnB3B7uTYj4dLc38HYynhBq/RrGjo39Qr4APm/E3MyxdZ
3jYBsp0cWlbgqqIsTlFmVc8ZT6IQR+Q7ffuvv3z2u5I2tthN+Q96XVSer1jIzOEl5TXrTo/+a/r8
+i0Acg2ebH1Mzw0ttPJNm0bCQ8EpVb9bg7zoRSsHjHuDMZ8YzxXdWOZVA+7ubXw0nfiewAhzpaxK
fJNmPWXEQQHL+mHEz/argKzw7QHc5MJTZyknIQ/FI+TShg/fcTp7XaYZ1ey7Lfw0p/8BHnByoIjq
1XnIB8eExWv9rWFpahLRtFU1ywCnscXHFQdztU/JSQQ32fgL54uoowYZtVAY6XdwW+PHM3f1Rzto
Us0FVv5i7bzqt1LBuDPo93o+H1ajOR4usVRSqqEIsW7Xka/0LmfXNhy0OaQYgGwpo7JBw90k958K
Fsxj2evGrEDuMwn6WSICfincTF3LPlBXwtRInrbIWp/Afb6uYK29nbqr/XJgNh3p5BCg92vUiYFF
cEzCkAWa+1cLas5U8xNWAvjcCp1+PcNJGGbLOUypAV8pgq8CGHvaixLJGnybUW5G2hcW6YSdM9Jn
ZY6k9CST5tT/x5tPN8yNXD2I3XNlz+c/XqWNutx3JLCNexXgxlHSPHJ0a5Os/5GaaZf1Me+o7w3g
ld2ktk69zbD24AR2WIwlc/ZVCKGWj15uBDnEHlRPtYHXnw36lZQEJ9vGHW2dfoDj33EX17swQrX6
rqjZYO9vAOe6jhprI1u6gi/iHKqFET1a7TFkjNna6R5jYkaMUBpr9mgDbmIslIFtPi+7MC3pcYnX
uFNTRTpQhOLJsHQikQig0WgIbVGrQpubl5tEYi+UcZxve8X5OPTFrxl8Ym6g1NJlsFudeT3rba8p
Xc02idIK2Subp8CgFVXraHA2C/dDoN/8REaC1lH7RBoobpfVB6mAJcwVhVsARrVbUzzX6ugHAZXU
MkD94kIwUoXuqskqaY69B6lzqxPcGYrpLmpXxpcPkgrJUtYQM9URnTanS4k28gKy1oJ2ogehdGHJ
y3NAZMnVJfAtoSgENeuxsGaNwOnlBSXzzYPaPSM3Jhl6aHxbEQHJmjm0s9cOkDhtziup4ofhWfQc
LEl7GUt6BUWqEXfSJt117fMqA2Q1SY9GxyD8gfsyyO8otqKILeiUxtGpotpehM0n6xFg7npT2TdT
xzC0WxfYVGTS+fd1KrvyI2wgtE6zcZdykglgBkk4CQ9pGBC28ByRWJ2ZlTYp38GlgvO39sOO9MY5
0m8sMe/RcgW9pxYTMFmXo50U5W6T/Lmm5yt05qOwrxhY177+duMlnhVoELjElpWd9FrTC6WmIGG7
Rk35uy/7L/avfOOQDY1Z1DuM/gp7j/gdXQnGTI56nPQ5/KPuXs1jtimBqcWNLhQDPmUbWBD/3Leb
uOLCX84Z3jdHXXAQFFB7ED8nmRnbrewGi069m5530YT+TG2J0etv2b5Cpfph/U4KqKPQZ/bStCzZ
jXKfkFgN4uNBAFUNFxwKOpxh59BX15aWapMkafSAHvVk1E7gkfppiqixo7S7WQbwknj1voCue2QZ
7TYovPUQyDwNE6OvHOfN9dEW8r8rf9RVpPAxgzlhKiG64IO8J6dN+kJnoM6FK8ye1AcSN0bTlJ/v
xow8P/s5lMOWgjHo1MqF/k1GKj1cxqiV9+SWXxqZUWw2XATc9jV5nUK69DOM263mamBFgFzLXv3L
tUYRM2IAyM/l5PifwmU4C/l39onqWYMpMkszdy1S4wNp0wQHoWPGwzuEy4aq5SO7K4dUNh7HFQb5
hjvLkKyE3UeP62HVRkiVX6uZAeKfagJwKop5UiUTc3F3cEZAjubVMcUGoby6becLYxMQfjQJIBfV
GlbC1wk9xv/PKUQLtmNYcjEXiZlo2Ro+pUmpyKFd8o8osZdxWw0ld3oYzvKb3qD7cJPnk3lVZ6LB
CHgirqZ3SyC7x4ao8xLCPp0NJ02yA6LZPQ8lXKTrGMTyBN2dYbbX317wKVHgUnXewIDnjuxU2gtq
Zs4qfcDx8jKWPhN1IRZYPQeorCceFg/OpArqFmu9W9W2WCFCrSntFRO+SOPGZjPD/P8HEUdaXs53
EFiCph/nc0XO6TTlH22OwvJGI+2+9FT8YwwxjSidvdIPb46tuaAgLSuezf+KJJlqsADDUHLCPA1A
/gR13GaexCcNzhBi33zhCodj5czoeS7msWwC3hRrmbGCAMfsRKtHBh1CutCNBrN96wlUNrncLajF
tLmKk2jPKVdmnKo2BY0Nxd0UYtvHq3FxdBuLTjoVoI74J8i2EOcHjzUQkq3nYNjrhYY+PskzNy5M
Tszj45joq6fneyFSuUDJekfCZJiShJRXyfStt0RteYWPmo6jxJSlqmdREW2QpAB4DV+lLca1VETg
A41XGEPp+nXS3F/sfHW9HX6u76SHW3UmNhRP9vEfklPMZ2bIMv0TE+V13+GmKI+c+0mXFCiZ+vla
g35Gs9CZJNDfqY5L2QSrw24hCxZwS9Fq+H2HIXDw2oeuYoImA1Rb005nsW6Hi1cfe7Q83XqlzviI
2IbHNF4METM9cYOLRseli1rfzkRd5sKQzdOr9XtQJzj2YYKaGFpiHH6WcY1DddpnRrK4dd4Apw3H
L3d4yCxl3rDqrdJIiP/cAZ8TSvqM0PLX4OWjaMs9MX9UGOjss79WPzc02qblxbdqlhIG+3LBr1E/
B4Y5hRKizvJAtfkq7JK/GOLMU5Ji7d523R8jhtfEB4AGTVDum470DKIAwi/rTfm6n37y49hTFS0D
AFuHU66wKSLDNQzLfqPNTuxv9B0D1CwA8jmYWwVvbUrQaz5/OceHm7AHs+8ubV4ysipr/dpng+pJ
syNgTtiTTAwUZtcd0qBYsnareVw1P+5mEheL2UuSRFBFC1DrYUvZOryf9Ancm5pNt4/Iyn4D7Pw6
+hnQW8/wEAEVm895AWfpfXplqdJzAGth8oCf1DgCnk1IoE3Owi7C2tV5yEmj+U+kGfN50caNHB4O
hKaKQ+KGci5FG3b8SiQ6y5a7fLWEks+qrzU1AF/OJfsokrLGkjaLX8LMk70OZjaHW3GEyxQoRgkB
ixw27fswHWpom6lx0KKR+XB8XRiIYYV+giwA1+IFUqFhE2vHX65ET7ulY9WpGAK7rMOirKxnv+N7
rWgOqZGZtBCVHVl2jGSO37CzPP8L7EdONh9okQfBXJVC2cPD/8PUnd+6KsDwkCOlewcQP831EAgW
XAN/d+RVxWphFYMG3cYuXkJnf3j5TD/NJZtA7AAIk0ZKf2TaaYP20ZNmV07Kv/kjlwzpQETmhp2Z
FJ5fiABarhTnj+HPGT+fFhmCd9j2JRekVhuIW/ge7K4L5LEfrFut5e1UXYyeYR6/4cmKLLD41ZU5
4mmmOLdj+bEJzenx2dxHI1aiIjY+4OB+3UVlI/e1OuXLJzTayVqGpAuiKq1Aemxy2zdYuHl+TLQU
NnaMDCHIngADqsl9WW+U9ava7H7JVvducviE4RH6XyZoMVZCIp9nlctmEd1yeI9PD03ACMCxSym3
AYvK3x3+G2XNCPenrApv+/KjOmqmqKd6vdfqxEwPGwfUV9RPWy6eNsfEE+pzWUyDTQllYiE4cPaJ
DCf2hTP2hACwEnEW1QErk/gZobYUdGyNT2rOiI/7YBUwZNNfGhX30M0B6VyXFv56uogf3k03m7kA
KqWCrOe699ewYxsNLYDoD8+YqEv2GXgSkez7VB5xdnvRM4TvfDsmfCSFg7PsSOP+tlH9A+6E1Ify
I4ntB5jfwF9NnZIuUGJpESsrzADAIFCKvar9amQaiY19GqRkrWWZov5mFdjFR0suHstFmxqmvi34
aCcq6+vGJzXLh9GZoDGWTXdbHeyzcs/a0rz7iXOMyFqlEDUPcDMorEzp8npWYXKRDXlNLqLlYLOe
nCg0IAGoep72hZpPzggQG02oty9UoiElEzOo9Pk2knbpPdvCJRTak4AUGBajtV2Q2N6yeejcreA/
xS2SYbD95gHKrMo9JknxCbG/6JBg1YpjTqc1oW/5tf68wSxb7yMK5VTmToM8WY/At//mz0OR4pdQ
KQ8TL9dvrlnzARUHO38nBj/OIHzNUOGdXjd/NrRstFHYs4rPvlH88lgUHefd5509g78PL6fUoM5L
onaX6ao5LggaNoqnn9Ut23C+AerH55AaHSj6U/ClIdg2Z1YufPliDApXTt8c5vgKm33jHbF+0OfC
6gMLFrKAQsRuV8n5NAWXFlv1G8pdd3avHelYjVxKlf882pvq5/vzA75HFSCCgAheJRhxNjaWOJmo
bvIv8AAZRBYuLcCY+fhvD89PcdiPS+CX7qPLUBxXRQdRs5T/maFTXsMYClbOuagbHz6Nk6hyuonJ
qy9+x9uoXsQcuL1Y4ItNZKIeGQmk3bTb8Ywd1MCG5/X0omEI9wnfooZxxYY8r7uvLrXcgD3RvwhX
eztiwMi5Q67ap5oEAaE5uk/QwE4h7Hz00efK9N3mgmGEbxiWBq0zhe3WlLY6OjXhahFJPRaFRF2H
A7zs7QuaVasbE/DRHDQGUVdV0UAYJKN79nbDowCORqv+BEFFUoXyCpsTz3LQ/z9osacVD6oOPE25
stZx/0R/4aQFNkrUHyLAP9PSIz+jmX1gS+HYdkoejI7sIGhA51iKNp9UGjfIhdGQQLDk27t3+/PV
A3I8Gf5JiGhp2TKSryBDIBh3EvijXTMlLEcDjNyaPsezUTvpd5KEM2JawckobscoCztCGEezhRR9
OCretN/lDgrNyQROUrwTstswQ97O9cGsETYKBa91vS/KqZpMS88F8A+g0ZPHFLPAlA2WFsL4ylJt
yyJ+WYupfqprcbhsADv8uGsQ/xvXhhZ5I82NGLBJ/OGa12k2psL2kwU6FsPbC+96pF3j+2nY9wE9
eRCXplFCoyqks0jDpX1It9OwyN6SB0M2uFDpEmIH8StzdSY7UfBcMMaE5CRL6H0bYB/TqDdzoHAP
fKZaL3GNPt/PPb38UIfYBEKrDTNrDVfsu9l1oocqAqRqLcm0vi1Ra7FPiNFDOOrIAT5ZmsCkpsbG
mJlKftyUTyle5eRPSiMryc8R8W46oiy8+YL5ADgYBYPuAuvjmIETGJj+eodmr0TIkJgM8HO+vQAI
/492++9hg6TE8y3zhvt+f1E4R2LjZZrFfaSDq+PfhTm59VDB9zGt/Hi2uzHl4GEvSJKlXuzArQMw
oh+i9rt74qKIYTH+Mi9KS4bRjbq5dfPcwhJjmshBgNNpng///Gftve2XLk4n4AadhL7XZlGiiXU7
aErs2axlUF2yN8aTuaMNgZUEPVWLMRR7tVDiumhEjNncrCNarDMO2yvb+dvKKxGVBVa08ArqQSrV
rqHN4eKJf7bb9qDUqPVzQJesZyOzDsQ7o7/1KghIGWbJ/dDjMHoCndmGDcLd85eecSKqm3AVoSXO
9ObhnYGbcUl7B14ATu8lvP9Yms72HLJMCChQstf3C0oZkEaRlS/viYZmq9spQsvQ9Kl8JWxqzsNW
xcpEazo3bDCMGQRutrr5vvI9IYtryllSwU4tj+I6r2xYSBz8nD0CoVtT06vJyWZuvjcVOAjWwV9v
siiH4VIkLK1HnWTywFY8As7BOgndfAYBpFemeEGj75Yo8JKROdgyX1SDmsvr14rGLSwHb7NSl8v/
epmLdQoLSc/97zmPx/tNMWiiWkVKy/OfhjakoPhLR9uX+Ws3CKWtZ4aiAMhTYKa+7p6l7B5OT+Ni
CFdR/moH7uhzwi1Lw8/kmV1kkiLcbf5InujB/rcJx88F26ez8EGd0GeGNtoSATe34FkNdyfaKiqi
BhvgawYJ86NegKi2ggIzySlNGPNCrQA9dUVRyNZmx5psbVkN0vKAlniZ2JUBPSi9Qn+cqPrbx7pg
M2otHrMWdkRpjUmS3RRz9yUMWlFHEKPTpvOjdqO/vROfQSWENLYDDzmlu/VlasbzYA4LlgtniHVO
7vxvyKciC8DJSiFMsO6DpN0t/lNXOoRDyDLVyziU6tsOg2q4HqHG1VLGqOsKk2nGt4+PxpUf5TIq
XOZ1uAuow0n9mOdEC52+9mGD9fuXnVxJ+jHf1fgiKYIiyM3LJxAABOi93X6jTof2Oqhs6TECvNW+
75iI0QfvMJJaDRuF0XtaU4fSvKYsZG4Y2Pi9YOu39tRXKRaQMR3lzIZcY305f1+YJVpbsuaEVsIu
WT1JhZrLovuJpC2HMIrJ0HihUCWJ30k3CwjWwxtBpGeE/AP0bwgVkF7eFwaQj+shfoEXvqUDs9AR
2zyVzzVKJuH4MVKpq7c2nbAKZHwfJbBzCL8ET7+wyQHest+Hj5ngAzC8Rjtu35DGXRpEiBvz9L34
lvcetOamVxRnFpQF/5Hiy9R4qSY7F4qXPcn4zDFOrim9LeJDm6qm7d23p1z3uT/56G501fppjlbU
TA+aqG9rzs2bx3sbMn4w5RwiO4OIuj2zbiVESH74ZBeOrlw4pFtJfPxc81xAhMh6qvu64silEXgU
TxfRqyLpnpUtJ43eS3FjoiDxwPk80XsVQmfxawzK5jMVrF/uIM/baS62XCURS4tjEWrukhZGXLSv
6Lw2OOpu581DRnLnDyf3/JyYByztDjCo6DDcsO4pF69BC12vOhFzckNvWRDN6biJcydPeho/vwMT
iikQjj6AFXVtouHGE1b31IEmvC98X2vVESRASsvz6uAGvlr2vhwcQOuXS5p3x1W8QaKWe9TuP+QT
QyMzxd5jbbv4FFZvZUQypxTx9c02juT7PTf0lswCBuEu7aTtvik/kymSmJuNxhpicR71zjwnZsz9
5vG3vE4OUSggZr5Y+4GPyb7cvKieZ7k9yNNor1MrN9BNYvmBu5/kxn3Zw98aQHuAK80DvxFTBsZm
O9Q1bqp7yFwG5qosAqT7aZo5CQQHR21TWjiNbXMB3GhBROmA3fepUuxsLvF7uYkWqJeeTBZxs9YT
YC10WcxtcZE8WZ99dI73c7vucbXG3IPPOTy///jL93XwfYBFBCbXqOgcCjtw5tleYOeKF4Vv8Io+
VHqqCKDozgtAxmLhMncglkbXYeg734pRG3kvDyLwzlYUuxlhTfKXMOhE8/a8FrIG4FSHWq1FI5dj
9QXRrYZhKYRJvwb7dGhdSP2pQ83Ap9GxFYH1KmDBc6YdSPdjFNyhuChnlwbOKfJgZ08vJkJXl8nx
B/k3ye8Hq/spYNW0Z4IfaN51K2B6wjVEkTXYN7Nf4n7Txs5ePKXaomxM6ufQK6wPXdfm6GvOzWif
5iqQOqhy4gV8O6c9RXg1BjpxI/+hfW8I6kDhi/TVyjTthGVlzE9G+Zyt89XS92sLw/rQiK0AGK3j
9blsnplfG/VNjTCQmUbb9aQpYK+W0i5Rvcu7HRDoX2IgY5poMNhTVbYtJspVgXFpSEtclo3t8jLK
OhWRt8UsQrFhmAvOS960CEZnz9FB80X1g3A76OEnFfIyFdKxLWW/h8dsc0JPnmHlt5Pa5ctFLzFi
ngrAuOV8dYYavMCe3p3MQmlXYFaXChQz+uyAFFK10BbkJ1l9fBDwllVUvT06Gi9FzqMRGPReINkd
6UmcII/CrIFIgRDXvFUqwDXNw+cVEoaUnjktAXjYd1xt5xHQ2hhSwliq0cpGwxgiFA5pb4zz5JdY
QBeHfECj2ZWmta7tqQvl9sGxd+0srzl7jymnc21BfT/HepjQsLucrBIUrhhykO22J+dogX/thX1o
ddXX5yc+5o84Wh/Zz+ZcraKUufxBilmG301YT/uJbHn1SFdDK18np26TQlZ+475un9XBZCS/Qhym
G2qLaa6Jvfj11n1Plws1qp9p90+u0fgMvXoguSRshYpc0WnwFenPQoiBI6vRrhKRfkVB18K9GbYh
RrCzU9asEwWMVEAgbhTPc+FBaJ1AiKCcZCHb6MTQ7crCd/X6PHELQPF05bzE1NHfLJH9U+hsGOJy
C+UmD2A9fLQrsI7vMFPlPzbg8tciATpStkzVuJjzsOo3mwiDSx3eRELhrS9xKrsplCNYUEopYYcD
RKJl14yvB7FwpP6gaLr1ucZrLfGRylrFuBm1cC6S10E4B82nhb7exDz+XU99RMWBczNve4+0FgTG
KxSlfUGyl32WpCa8MJlLk5FVPO2rjPa3Hv0cMcf/mPDiys4k0XgKNpBghZo73SGeiRDrh40ma7AA
6dZlqUPjAhe1ED5znyfQSm/7zfdzIZHml4BnW3CwCAxtQmXqqNZxEVg0kNwnLAEHyKO9W7wMobCz
xySHl//8IfMuYY5asVUdLzhBaqSJbn5FCp4iLduC6La1wu46xdK4/5GV0jNXuYNtoyj4Syx5mznz
PXFk82n2AUt3XcukbG2jwsgx2L0Ja1at4fmU0e/m4U9LVbu3fFYtIrVXjdIRMbVqx0LDWBy6HRdf
p/hhrxcG1Yh/AY+B9qKfpFchGlFQ5dyZ1cbHJzcru6OLN0oSVWppUxYy7h/z2UXw+XrYdaXqczRP
Wf4N0Wls8NJSEwA7yJU1/c4CtdSWrJ54fVeUeazxAxQrgyCG0QOUq+fgW/L9w7k36VUvygdLRPBT
bdTS9jP3lGsFC4j+kooPF3HKjMlEn8ufXLvEjRfBQ7+i0Mv1GEQcTDhzkroJ7vhb0hurk1VFFVIX
J2ksRtiqmXG8IIit0w1CRNfBT4JLBtJJlDwtz+iZ2xuaxBGdGE1MQchFLzcUAsh9s/Ha6nAHy7BE
bnBKB4OexBUzlfheoMZ3mmVsBFtbc7ZPv6P1insM1YRhSBHQUtLAgGQRHAehBMibWCuqDHcdbH3O
o0wwNTU6Xw/9zp1ku0tEq8/dHmxFF6zmBPsKlMs1yI4g2qHuZgS+e6aLHTwBM4gU4kM7FTTq+BhJ
H1hG/lExuJyItaXUReFHPpi+2hnbEAuqS5A4VXy2JX/ceQCgqftqU9lwbBmYRQEP/TV9oUHa4VyI
SEHAlOiGbaN9ppu1yPuRffWVOhLy6Ztd4KAe7Vbw/SZMHyeb+o3e3VallZHj3nr/RUrWjt28uE13
wW7woO5R9dS57GSOVhjG6AmLqcOhhpUBm2ZwgfL3EvAx1fh2g/+33wnYg47ojFu9q7WbO6ufWx1E
kA8TD/qEMOhlm6OaQsdQMqw2h3+vcq4BO3pQVCTKCnZVidMNWS/eP7asCGZX4S8GGSMFjsGvsJgH
5LC3FWpmkrqEtqtYYHaiIXZCEPyqoVwBnsUz1LTHMJdZMakdWNyH3+M4LWlsi9GEWU/2lNq7Zd8n
2v9fBFeWYTn5cxYK45jm6AknP7JVfNmgzyvXsfFH0/571PLpE/EvCqt9kFXZqkI4PT5QrqFW3Aa9
SqM8CcdzPKbwe03Y7wPxuF7YzxG/a1fKhaSQxqgXqFcRKoInBdU2Kg8Edyfzx+niM0tJH/vQj2s3
Pq1gaLETJajZzSlDqq0T5wSqM7CS4+TaynOS3cDoM2JpRmvh3f/qfqWDYwWdzE0N9Fw38NCew9ZR
/p/Pnh2VyExxRkAiPpAYR/uNoKCC5+u+GiSJXpn6hij1czOquI+rDaSt5k58RCUGu6ND3ngJUU/D
OrIfJTEOOv+2Oh2Z3LbjjG2RllhTZhyrpB6FNZDG86faOfSk6mKrKVYsz7H6SoIGKHBsZgABOBAH
SfbcTIEhxkl00U0gCkusocexigKaUmSt9X9wMtCtcQ34/uonMVwzUy2qb3tnynwN7sGgQiwVTcV+
jj66+clEd+ILCk5xn+RAJp/ZzyyGrX/n8LcAb+k0zBEWyBs7/Rj4lTlSG0B99g1KW1qPkKPqpXfP
cdgVYaKfsmeRGWSVMOx3Yq8t+In/6w+93buoCBRlqwdrLKjJwZyB40iLNMLjXlWaQvpxFIGYUsaa
YLK3G3/jfGwAlUMx9AAhUk35190R+C29VHe4wDdWO4kcLlXRoh6/CoIPvov7oxRTDsHxM3spb84F
ZDCEOrVoKQ6oYKQEdPL8D9Z6ja/YlJmBmlpkph9rBLs2ZIfq4udeE488Gt+qRCiQp8ixI1sUFDMn
/XpelDwy4IgO2hHtZ9NPEmrFxba7J/eQkdfZaCCvwon3iCzL7LRuo8E8QqHilkFA7+NIMHcVXnyq
B3TSRmFQiFgDjxSyM/J+YVC8aRVdS3LWLI9pChJVw56TBmNfxOrPQbmVWb8wKOJP6wMFzLEDGTBq
jHoLJbQtoMH/6ylNAIcBXu86zu49N+fTlPRK5auGk4QR7TJM6YN2Tt9pgAvFZ9MLtvozuNKyxyZ2
pTfNRiaQIn7JlRInfzdsLViWvOodiTs2/zTxBTyz1xECvKTlYodhA0L3zEhKt5NpxehsaEUn7ESU
0kaBJhe1+eEoFwdzChpFBLiQ12xIQCt5yDsNVq5B9EkDX6NIiY8/znW0e27Om+btFGvxYKEUOj5s
0+31TKzr1d4I64YJPnix81L1lfUWNGmpBESLjwGW4HQwCTFBXCRdSqf8F/QbTRCXprQxle+1DN7U
AoUjyUm+seqpQ6kSRQdEd1PGstV1s3/kuEIhiaHJkBLYIJoRBTOaQeqSwjZpSPIixGEqhngkfrm+
117H0APLtp5/7AUy4cVfd6z/fTKAO+PUe3Yk9V5BKjHm0EK6pNW9bh2oRe7ZT1Zknsu0rl2zrQ4x
qtl3GWltkyOvMIKFD0qk9emXBgTOvXJ3JJdcWA7LNBz60kWC7eT13X6yJXc3p4P0cGkBXQukdFU6
p4ImwyMIozeQTepzc02nu2rIv/GWHcn5mThqJ2+fqAwGB9lgbkV04TumuGHHu2fK5/rGUMhGeHJi
yN22tEhstW7XTQul0EOKBq1drcn9GgcUNBkX4jMK1h96NLJlNT03MQr52F6fc9B5OE2XkpdL89rq
2d4k2iPYmnLMUXbqJEsQ16ErsuyPdFnH8fm9SdN7S7+U1Pivh6PIOuTo5BDCRZQ5ZLk6leoi8Pkd
z8h6vPbsaHLkKooTxo40Jm9+jUJP902AMMWGtgz57+487vvSI5FE7qmW5FaDIarhsxEk5MJdeQdv
t+uU8/kuk+/hcQbhi0iLDGmJoFcrjUkTqU3Ccn36qwuD4XgeF6NPb4KMNltxpeDoOxQjsNET7uN3
Ey28O13mG1w/leEJtSxO25YzwqIuVLZK35zyYq3QlNl5ujNMkleM7RLY1KIshkTU6PHSWHmb/u99
U+cvhViXOoDOOnZwfuFkXx8EzBTepyun/AZ158yA8CKPuNQGccfLLUw40plCQ6gGo0BHP4ffEWus
QPCJH8uJCP7y3Avso8/qIE2BZE+Pqk+ZNjVnRJKkWGtM6I9gHGpbM532kAYSRbhHPF/Z1ZhBwVCZ
dx2KfEOyg4wCqMOGQ6hty4tFW0dUF9bqrtabwB5wdO7ArlgrPjnywXUhqVXzYcm7aE7SzSioVfKh
cNiMwpDg+cDW9cy8uvULUb3a19Ju1OjBbx4LhK8IAtW/fh0WFFzNUI2denk3tGMLR/mhYJpVzULn
NfzwArqAvRpITjGvke9sfHDpmOxGWaKsv/wedXzgrmu4dGj+yKqS3Bi/z665rChzAioBZji4gciX
FR1YH0EMzlKnp7kluBmXoHZhM6Lh8UI8no7buvWLrGQym9lwVV6PIC6nAEol+Gpk4PaUASBRhMzN
gef/VuYxiEvxH77iQX55h+4WQS27tqYzLXyjSonSLSZLwTRF8IMVfoKbZ3atjCqCVsP/PwTC0vJ6
p1Qhiv1wWPy4v+RUDQ5GUHfNBxZ/Ai0okYCjt8BREXgyk0Vw93mn0VWGuw7x0I9QJri/m+C2De31
VDYFNiq+xKgXx+3rK4tL0YlBHGHmaJlCifU182549FDZBJ5B4azz/BMaryYLDd8WDJEsxca31DdP
QKbiYSD6aKESIp8zQEDKWVvlTTahlqUgt9nALuI6Ana/tSrxKuykHjJnC0RsaR9D8l+kSRXbnuLk
vXCpUWO76nL+SUeYy1E8Kr7rPkwofcL0Ej6k+Se9LVNPOn/sdCXdX9v3qjgmYt/KmB4KVRn5Gf+8
kWD6GqBHpbqfXZIWtiXf5pru9alCcgDnsK/HGB0Xwlc2giGutE+yUgYbsgWVDQH63Xn314cEjjpv
L9nDPqN+xpS62F4OGUue7lUGWkbUOY3DsjdJ+/i062Rgz7UU7A1tpw9GYfH4IS5h/HQN8uSoNFgJ
E4pSQyWg7Vrn91zeFZywlmU3QjCLh6kfKAP9ukMVPWVoAgF6ixLhcwmETxMF3q6QFaEFrBYcVAwr
JXORz/iZ6LpazFn8tlitO1MVxoJNSg2l08/ATBGSjNehtWfeODFKahS3KCfigIctekHXnP59Oxto
zKC45YPo1YpvbgmR9Zw4jYBVfqGFKmHyRX0QnyFaLQJpE6guAWtwOI013hGfNV9T3cLSUmX8i1U2
ouII12Rnw75w5bX4oRaSYhjkXYZ/qAai9gE+nVMb3SskHRBKrvK7y4vQl1bV7JY59gNxVruWOQWJ
soP3y53yrBh7siIjCw9EalznP41u2PAFZDTKhzgF31iGx8CEVB8uoZ8Q6LO1/4uVDYoRNas5lQjQ
P6l09KB4rP2SSLmnkoeqy3DaPPxMwtcKXVkNJRNsoxtSfqz2te2HnsuC910WPs+sh4en6OfE0esU
RwT3qs0iudy5CcJRpuEDy84nxfq/L2Yz4G3NVCB5xVDAWnJX2vRngnSBtVUpUzMRNtMSJdNkBOyR
6xtJDcR8cqB6FWNCwcJLglWdRG/56z7h9JgN1NA3UpN5V9KPorD6/Xua+UBKJBKDU4LDRTwIGgAG
OmRAs1Xx1uzeG4RH7xh2Pvjq0Vfg80fBI/SCFA2NTz4PeYjCAS//b4bj4rsn2beMZejQPczS0Dhq
viMOeND2vtauv0aPo4lECrwiV9nNqr+hNbKPXBcCHZe66dwYZmeL0npMJd2ObWoRBRk2/cXOgUQj
MYwch2icfGthkU228UPHaw5E9YDU/E3WrgtAETDCGUuqV6yfbxtKzq1QEGWSOW6ZG2zbO4eGF8W/
1BW+/afBEvf1V35MGAjml4c6+Bj0kfZGOjzYwuI2+B1+wH/AeXlc2fDG3ZJLYufRLCHk2Y4LCNZx
sKKfgPW2qNwThDuIENo2cj0A737MRmSgVCb04OJXngRSbZ5awLTf49FxbkEJZiRGMx45Cc2WU8pH
axKOgNs5XFEP972ujZ6VHaZtnRBnH5eWd7KGg8X/CsIQaDWgSGGrqpXiJ7q9SMoLOfUTNnWce6k/
kH0rL2nnRlv/fCpbiBCybUUMzpKHsK0VwqgL/sJpflwUoA4c0klJJer0asFwoPqXQ5QVVyjMN5mR
eKPNM46/WHGuuZrlaOfD7VOkl6iVxFk5zwcBWDICH7tLQcUhTzAralCNEGINwCZq7osoissk2To3
whe1UMRWPe5LwEuHcREWQ6fxxcXmgJouJW4n7XO+weAV8/3gVRKgKosZwBjggt6NkQjyYJGjIQXw
7JtWlOWxi7rfupu1wNl5YjEvIbvTgh9VDQtLIiCuX8ffS1RTJBPwXKRdEVZg1lE5OenKo+VCdrxP
GS/rJ98oay+0rHKX4E3JwIAIm6tAS6K4qs1FJaiSdcPIzVbM5Ols/Df06sFv2DdHgmDmiYm4o0nW
s6Av0mmFZrDrm7LrU3e570XpV7nSqRETNpIhmZio+c1bUcL/mT+EPNG5MbZ/p0QQ/ATV8FWRA8zL
C1uKSRPdYwPP5YSVJtgJZo/Nd55SMhA9/j6qsh5C5Y7P+A4nnA8vX5COquOlTvmGYg2Mgmpn1oCL
X9dQ1uv2xznaL0VxS0KeIV8mGDpaPKrCQWir1JKB2v8eRL9Qd/fFqI+Cy/wlWiYj0YTUYi6a77uW
chJlrVrmVODpHRdzPDn8t3R4vZkrCZ3S/N6YEKnLdwjWU1tc5aTiz25eKr1Oc9XMzrahp/VodKI9
c91MDsVQqXH/twtir1Wv/48mVd2fH0Xq9HS3nzte2V2DQskMWDQ7mMLi/5vKCdfDMdRn2O9sMJWo
2HWV8aTDA8E+QpoVhlKU8hnRHOe3wRIgjD6Xwun/PE8dyxJLSR4sAXsSxZ4cwCoqrADUQTLBI580
xYQVoUxgdDWwL0GgvJelOo/EcU6jKGVCCTNG/rkAFcOCHpWAes7EucSrJxIdLPUg2yghKCNzFWnA
CTDkf57DNZYKSv45bMQ0IeskPZYAj89xpROLCwhLlc94bU9lhYBjEeXtboQCeSuB6TQTNOpBVZfh
hbKFSVXCsPQlasDhRCeJPiB9j2gCPTMewe70K0on82Z9x1Uo/ybE8Nd/1zGajxBPLxuAIUoMnyXW
+5YrrOTJSJ/IpBto/WrGIppt3aoGn7pvtWkYiTSFiuf0vze5knfjk5KJHSAgD8PbyhbppZ9RF1b5
liZ3kkI3TCGRKk3nAWZX5McVKN/BvzYYGJhNLkUzJfkcp6jWr4WU8IK6b4qioTUh2Jwx+pmm+iK0
EPw1bm3JQ/Wx4T2Rs7/Gx5/lbHzy8I6AjHk11rGztgAYCafOGkA4aet8G7NtvX7OY0iB5NvlB4G0
vXIDWlt89K4G/q/bZxIyXJUfBUFAAsELjxkOaNAb7gY9nXlf+c5vgilFhBpwJ/TU0ISYac4ciIsu
AxLfX+9qfx5KRMWtOaaH2zvLlbondOOoZ/HRNP1kFKhDmyZX+1YlVXPCWu3/ovtQNFb4xDuo/VRU
XlbLfrzPa+WQoWatH5GuGcCqU8dYcUziL89P/nM8piKo+uD1cCZH1QdvTxT1PF3dMoetugR8XekH
kEInMaqI3LeA6U3sWK6ZVVYPS1Wl53sCmRxPg1nkRi/c2p5YN2FqXvb+BjPW1E+kyPAx8PDA4Ljt
B7tlmAir1i45zc96iRkwKQAZLtw/DhJ7jiL9YFWcrQco40eDzUEgiDASsofvPaCzrQIJxljHtV9G
adTNbtswwN99A8EhlNoVMV19BVmu0QIPzN5Hl3imMJJHQWsnFKjWLKjEiw597bBhHiSFmb3dmgCc
Cc7+3HJ1FtcRiPOTaaNRZqM7OnlZV7V+9wYLbnLpl11E89uuU6Ig0XZUmSkaspExExIf4EnWeWmw
REQKsZEZ9IGyC3mbzeILiDzHucDS7qpfHgyU4QxlRqK7Yy/kPPOjhLBKR9XKxAs/uLpVfNlNqm5F
NlEUS9GMOTDsEDw7LXmb+NCd63ceuNiI/t4z/4QanZRZdgjNJLPOr4e2C+MC2Nd9dRphkkn35kt8
UyYbpb/BEmmih7jDmFbr+QKY3OFfz4cvPeVybPbfFVBtkQGGz0gZX3aA1tdpIDuNVOpTvurx+b+M
MYDpml061NdIrW+NfQ1f1RY+DLQ7/Dv+UeE+jmi8NKK9JvrdTUEw+XlCSzj54VjOT3oC2GIeLRxF
ciI6C+u/qgZNXISRykbX9e1SO6rPQhKQZ8g0dBC1eIox07aA/FF+Zq7eUhLh5cDt8a+sKhLQZN4s
eqmDdkl1oE8lDMpWcgT7CObpz0Ul34y8vlfozd+mY/0m6nqwE8oLZcMxDrTyGuqWWvp2I99OXCuB
3WddnTlx8YZbBZqXWL8zSIVDi7+sdVYb9wP+3u1GtKdN+HAYB6HJde4mH/3FjtSKXW55hr9IBQUU
NrMR4f03Xbc4ptEV6YH5ibKEkqkRGeHNZmV8fu8jtFQdthEV3IQK0TKVHTIl5q1KptmWNjQsG7fI
R9YbLVPMXW3peCodNBFNQEw5yxtXnAsgTOHfh9UskVjUtRTzCbSqK2tUhH6TqUAFQh0JMMbJhF5g
+68svHutokU8EGd2nEppgVuU1+Am3Adu1pUSIy6JD8xnU92+LKnSIMHWUB+q6FTbhPHl0C0zlSRz
LW4WAPgzT3FExukI1UvzylAHs3pRCQx64PgkGFlFTqDdrVe74rjEMHfDh/k9nEWuy6LNbpADImTL
HtHpwJrv/nUxBShxIT1TCsRd1Ojax7bfv2EhDJPHWX29yikckUMokO0tKqsCAZ6na3kJWwqe6zNr
zmbF1vze0FuBt2RAeekS6fbBRXBrql2HNSUIyF/RyfBX1Eqfx8zJrG51TiM+Ernw1LAQDC7aiwx/
iqY4UL/gauufw7ZxkIrJmrHxko14yFytzhqy+AdIFZSh+My72+se+6KcvonxnqopArcDH+VbN66D
ZLB0wBwvZupUd1KKwoUfEn+S8e9rvC9rQjtCp6KA8Vr3EtbIPquDTcg7w+P0q4R0YA25Buw3tuDD
YboL10BZPRrjKWYl/X4SD8tBteQlSCjKxIi8svV3PctLot5VK9Xo3JFw7bKLwL4GWBCjGMqec7PB
tbB96vY/m4EB9X9lXXdsRJYL6DS5hi6TU+xEjBVeQ9dm+Ts+vgaED14yRfD+7+5l7CzMILuiXEDV
NxEFIoD2HOJ2FRrg5wuhl6V+kMWcPgU30olRvr6RzPy5uzYRlK0GE+eTm3FL73Z7OzTWYJybq+GZ
BkmcNzG0I9KjYVmCuX6hoXIRae7f00m8O6zPNcND0CLDFeZRn6FiDWBKEFMQCaBzBokJTwrnTxHZ
HKpWECgi+NqkqYlcQuQTcAsf2XOgPmcWifFs3Kel2rlJJQFVnKq1EsqLW4knVFbjyZdwD2pcRei4
XWzQWBNnHtlo1MRAnFRhBxlvbk/cCGnf5Th5XJHojuwIFM5VaIHNU764t3g/haT6wchoIxYrXXKa
XFXzSVAegQTvGUMtdmztvVdgnpvzVUqiI/qJvXhJrHVpq4CsQ4rbHuhN3rRKQm8U59NaK4VNBmXd
dvF6gVYkfP2yyMLFKTPT6Bu62I2uTc0Bf2ztCFUvw1p1umF9rVsTfCVUeeNlGW+dxA3oIsWmYset
oOc6qWd46CrSLlimWhClSca0h0q2vQn1Dw8fsd6ZtsD7YIjuW8+RD6QEzlx53vG37FunL9pwbBuq
LSDF9Ca0jO7GcKxB/svHlMXTVjeae0orKNbhxHiIXB5DFgazVx8kalXGxxZ48iLxyFdPehC2c0Eo
MPdwdwSHJqkpnXhTlzZxVPRYYGsU4KoHGqqju6ghLN3mD+VS7R7gl0aVMKNQ8d7+e5jpsd54xH51
rJiZ8C3Ix8UWz1UeZaY9BZj8iQRXDs0VP3YC4VE6AEpFNQ7DBUsH6afID4i0zD1sBRv5A5IptE0v
zQHtNH77vtTK4jv0rD4J36zyra0945C2wch9053Zmpiw5BHJUS75g8DuI9VbHe6ESXG13Rpjn8sW
TlMeTT9meXHIY4jsMCfR0a99J2pPjHzR64cP2Hn6Zqlc11ALF159r89LIrRZ4w5znu//DR4r9Nhy
18wJQig2DP6owkCROGTx2O/ZlpYkkj0FPJvfoSw0lrgmHCVCT27k5Ayoja+WnG0W4dpLn6xfGgWw
53St3GJr9o3C+qK2QCcXlJt/4i3t/IDNJnnxjrJp9N3GbDIqZqVQK1N/mQ7rfkP1tKzDqSDWY6+/
5dXksLita/jYMuWxrTPE+elNIBg2BpPI49pxfRMIfSc53gwCzn6xk/U8xrePvE943BUQyhkXJFKG
iMQQbS3EBIu7llTLAN4DQSrrkB89NH0qkbLrVNsV7XStQ73cvI9FOx+V6/QMLtdPEUK8/tp1bFnJ
z8VLTKncNmS+7wgnhzLvJ/ZNb2bbGZiIyB+KmSguSy+iMYqwgGr4ZRzaolW8FD/xtZaA4oYqcfyp
iwLL+GM4lLOm6DMEeweY8cXvPxTbgShLp+7K2yOCfMPv/cDlPlr066X0D88VHrcAuqGFYQ2FAFxs
NhLPKZwYcDTsA+Jx2W7E9vJVIknSmZvR92VLD/g2QprhnJlfzTjCk6T1ban+61uBugWAG7Oq4cGC
QUXJnIYoR8OMntkY81SEPag3EYh2GdESCOB7yFLb/uVsvgVNKuZMImEVhmqYu823O9WcEkhT7m4w
u6FI2syPWgbtzlMyfR+Pb8KW2aZ4jcGh9xSgmaaiAckL4YkCnH/uPmD1H0pSUGOJTVa9aRnaoE5C
IScFf0bpj0UytaHxK4N9waxVRbWtnEugjWSyQ1cxpXsQ+EQZxDgHSjpnnntUEeJcRQmr3Zsnv9dT
tV0H2PmVP8vvApG7BE2rE0iY3/TKxWwgvbzLTgNs8yPv515V9QsjaD7kGF010nInG3o8Bk6nzb8S
06mbTw7cbOcWCjcFX7MHyxuytKPeJDg3AvvP/cOINTuzD3Jl8jYkWaOYNGj6tWoxvCMlmOTahaUh
OJrXkSJLFS2s48mShDTSzA7zOIM1SzAH0CM9ccD2KiLzPNeQWpQS4PqYQH8GYUb3Il7QDBBQz9xv
UFo2jQZLl6+oHP6iTdwqEbLBinz0SOByInZPvoRLHRjZjAQRU32EKMgh9/f6D9SPC/1TimPDmt47
29B8MY64876xzW9Job6G4S3y4BmkXepZ5d6+/qyEA83Vy8fOwDYTIuR+0b2kT83w4Q2ThhSLdTb0
3RWykrjen7u9PiXenxxcjW2s+XZOKDu0IqiX5PZscGMgmc4OOwGO2VJf6Pt+hZGInh2JFBbWC9vA
ZxOOzmuPYfpiNAu+v6tFgtJamrbEMh0YpjpMjZMDQY75oVnbqx6YZVzjPYZxYou3HbgZbsblJjsW
eHWPHkmUCheW0KVC+PV0FpReJj2iBpSQSVu2xqLS6TJoHOoB7HWpeHrPYHEzbZ+UoJvurPCOfJd8
u3gHr2sSG7FJc2E0PLMiHwWgo9sVUX9WPKHGL4ryjLLuPeRauU7PLr/aSzDx0FDSGlXNe7uC6COf
EFlJd2MtSZvSrZfy88ChLW+EvxNDVUj8z7fcnv9MyyxhQuFAbciVMTMjZtbWOb+1+vUp2ExMn0mR
oouId5Iw7dOZciTxB/lZmjSTGxif134+GtZcIlRLsq3BnncffZNdj4gOkYJiaZ3UN9e9pPRYV3D3
OOlDHoxmneBZURqv9wp4F0+PSrcA0Q/i9lMYd9eCh4O4C9jGQMGrI0eLGo08vWySTvLbFK9AZgBi
+X6P3ikeOshU70anNCoaRWFfDUDuGqgogaPGQ2OKLVBAzGuThAVblxsKaD0G49qyZntJG+nxDkFW
saoHpnauOS2SvIr/i6yEXVqgPbjdHOjPkTeYU4Do5e3thnvEulZbpGSRA5hVH+1a89X0gyMKDFzr
TOiN7+0jmHf3agwrj81dkyAhA+jn4r3hDLlre0Vj3kSC4uzhrIONUvuBA3LU4KC90gWMUdu4LHKO
gmc2+cH4QTUKcLkrQnjfzRJkX0P1cxo137SVeV5krIqFycxziN6QWvkvm9iAOeEgWQ6tLKCynNpp
9ebJS9xFVpR8AKtAEJIpMVNqUEnaCpchfMkmghFsefCCZNqLhzC1qqHMRjg4vnk6RZTGjTFHivpm
mXRo/6hYvC7gBQ3R6Bf9Ofo65eBbLtQGA8bpOFXDbGwZiqX0gw8LleTxDR6q8Os1YpI3TcLOWJut
nquVEt8nB07Mvjbrzq6IePg+HtPmHeDJW6GRvHiUYsA7BMch3DPeVq02UO4ytqOySsxK+LbwdrpM
kVh5WJiGHsrT0a/H/PgMrhC1U8NCh2xTHdaezBeCBg/tq1sswYcoGsMpuyI3BneCA7Dmsx8Oluml
bo6jZgAMKu5CF87qxtLGHunKd+eUXWlb6bMeRAkv6JjML7hUcjQD9So5+LfeRFMZBx+nc7BAlMBI
I4RixlXBrXbzu3Lp4WrRrF7A36bFHQhHzoA/LaMN4jYxpp6NPNRLbwXV0i+7qUvRipOl0GrCwRwt
5oq5mG8kRLRK67hqXUjI6l38LtdDKse26HV0Ls/XS54g0JXtEytYmuvkbCxRNCa0+AIhEn/5jkiS
7Lj0w7DzVKE32cl6Dnfipu/wfCLyigWGyV2hgmXnfHzo6AgPURlIdyQKOlMHS04Gl8ZSsrmYmXJm
Q+nLh73L3wP2qnms/DcfK+jlKtEksnscApQL2Ztv8SFWIpB8QZEvg9kY61yd6TsDMuSgdUBUvnyo
TD38t7gnagdYFbTDw7vGCS32ZILcj2PVdkp+9WlNyOSmF7yPNGNcZ7LfaJJcvdaLR2W5tYQlaSso
vzNEhAKsNhUiC7NbEGLZbKpXxePL88lWvxsCoAfP3EQcXDxh8u6iwUyZTMuERJYmf+pMDLAgqA6L
y4ODWfEjadvGBjEZTRFZ6oqdmcyKa/NcqSFO6vSPYO5zy1IYbUbTv206ezYXf7JfmMp9/PTEjKvq
avnBUfY0VevKe/9e8TyxFrKf558wuS52Km1oeehJr+Z/dGrKLKzhzjsMDk0uKQrIgmfMI+MzwJfz
NPRD+YUArgre5I/1KP0GG/xkFp/OnlzggMa/CGnbsGQ1OQVgw59AJJDNpvBkp2C6o09kwka3XHvO
faBe13MGTsPZQTmEyjSFVcLL0GZfQ6r9eAbWZTmH1Nrur5QZE1PW1GVZyb2OspIhxXflg7fYPSde
KBYlW/UBqo+38ICF4R0wYkp+I2HwKcNe+yLZjhBHWR5wOyihhmCPYIYQC/PTAW9jiNkPmIYFQNwj
+UXbxWaEWcqd2+AsI51oMTRaVaVIFEEKbFG510aQr34j6hcMMWTAwMxeNjrBudvTofLGqu6YtVCI
Fiq6A+OFUmhk0ceNsDUXlWSRSKn/+i4f5VZ7STuunnWg2j0S86QOV3RsF/6h+hYCXSBhCXtiur6x
0/oXrIHXm0pE5c2c7VfDNChEPGi7V2LqNYHPe+37BLl+6DopG9u+ZUxAsarj4yOQt+aSH0olgzXX
ke3xaoNDLHXtS9310bnSNtOvRykJqAsKuuMjndEgL8+w1FEjsV1+cXKhYZtwsEshF0axdoJT+z+l
AUGfATUtTw2I7JBFP/mUL3GnPZqSWZpxK3e/YIXKN+fjPrWvY3ZRuuUMvtZtHRPfWPvwUvrZ2oGl
grlOXpPt6rs0B3cZqxyVaB89nX82C5Z2S8HcQ3ehiwC+qzZ7KCCdeVxL75XDAjT323Wn3xYwsD+L
XXGAl1eoNDd3YAvpSJk24/VdSOCdUUQxZ2YGC5ByV3g4f5wzU9+f2rbndCXDCdQxkD8P+tl1anL/
wmZkAhqxyVGAeeM2BolqAHMWwo2eKvauDG+WSquSG18nmYuaOIn3QZ+ZAkFZDee5HIOt9biKm/QX
vIfV9tadRaFNzH7+PVfAmc+GCylHrXygatAPQ2AAv7ui0VCTJWevGAStchnOX3eXrnZvO8sTKuKa
TDRpJF0SXGbiNZW/3+w78GoEhZ5vioKOApU+2Z3FMvQl0JGo/AdnB429QQRY1+JU5Axe1iqujLfr
3LCwuxITnsze23LizbR9sa1YiV2Wd+AnQKoW+BdmUiyzjSDfdyhEa22QsBM78oVO8A2Ay3oQ0hoA
mDEp/StiyhSkIqCAbP3uZvJzbvevNLBfOEmtax7SNKcSffNuG3bhGRKDooJkDiYw+cWRWHKnwx/Q
O1ui3iUaxcE/S2RbkXw4VA6VD6pJUMTpp9u8VvO3uWYEB6BBmvKfQHdixliMQK6TDuEXKXcBRlFV
fwy24nWaA+9TbTHYMWD3riBts3Q/U2qYp1YUFYaHgYUaBINXoxUJodm1cE1bFrzmfsSw0Y9a47N4
MLTJkM+rh5elTcY3GY9Ghmr3Uo4QuNjCRsMoxzQVX9PWxHmA5pcE1hOjyBkx0eOqX1k1I9eKLhj/
Fy/fP/K8bgfYxFISOYrnqtt+tReSTGuIjRMLFnwK+t1f5ar7bfPKmvKcGjj1uH85ezrJV9XBY9My
vZ9TMFyWkzxu+qHTJT/6udv0PL5GmPJDtE5fBommGPlmeLYOe/wH2eI50Eb/sogw9ObnVeEbWBuK
k6vexzrcRGVLrKyDgbdoS6nsUGFXu0nu3IGT0qkpT5N1ewbkMmB1ZDOtzmSvxn8DB0m7sS4oupAH
eGXHuVWb/uTSwzSRdaOKU29vHnXQ3HuH97yUDsNqEU6c+qdF14hbL34hSgTsWkoZhsWEFfzhoMzG
q970zf8HZnvwDSZLbULpqRkOpuwHPR2LDnrafSRkW42u04DsrUwRCJgG0V2g+TJaWM17ZxEglXal
la+7748bFaYZqM/NuWzOxdOW3bZZG6MsofmM3TqzlRbbW28jc/fz0iE50Gkp9yxGDCfCsV9vdO6c
OadpniTDKX4wrx9B3fC7gmwpogi5BSiTEqmIqMrSe2tmtfr6eDdY+Lpk11ncL/tQY5ov74FoeIN+
YgIQ5NqdzGtk1fIeFA3dDM7WbuwsXpo+LxAgbWBTxCX6hKvkemr6ZJQZFXDVhjDU84+jYowIZK4t
bEMwqUxIE3q+ea0cPBF65ac1FhD20iIbPAPN9a2roqOQHeau7XFYXNiVPhGt6trquQ570snTsm72
4jptJ/S4kwpQaifVi6qUu72qWfsI8C/U07SOmeNsN4k/J989rHPitOUlgP1aHRQFM98WTzlUjMVF
9H6sWzGxLPytWZ3HbYhHjKrbdQcIK6ztQjfrwnkZONhlWgztlivsOqQcelpCUZnktZ9GI5a+/jAj
SRxGl5JFyr6BcqFUrmJcmkjNupk5FH3PissVWIUTzQZ9JQAmOKmZttGH/vkU+XWO6b3BybjkfDp5
a0tzD4Uo4PQeERFsZXOD22q/wPji95Xfij3F/OxbGX2mvX0Y/gA6sOKNk6dJHleWq17opIapFXI6
nm8z7pcNXSdTMSPten8mrv2/5sADJ92kt6IyoQX5eTff/OPO/mbtbDvyOTK1z+DOWqWi3QpzqXWQ
66ZNPf/g27j8u5eO5C99UNVwaq+DTuUEP3buDwKSIH2gB1bH+5U5RnCjz/9hjwEoqR8fYzy7RF9R
Yem+v0l4610jKg8K1Rtj7t84OapK07xSPqAMccpzrVqX1tCs5NUbccMZ9LVbl/yBuID+EQLz1R9N
jEiGtLy4BZlXVfrFVqx9k7nhuU3xrd0ZZ9HeTEvLXdeJP6n2gU/3fi+Dh+hj62thyOrFzCSXOCd1
J0Sh1luEK/I7/9qFZQx54Vi1Dk7FE3cTqKT8uCc1y8GzLhMHoT0J38TEdn+vQbMH8cuxeEXSBvMm
CsMGm54u82GWLtWpZSproB8z+wPyjM5V8wRUgCRZ3BeQyIuk9lY2ZG5/S+Tif1o5a/EadB6l0tz/
W7T/v6NSlKuMy/pKLGkiyvwTUi5dJjet0LWN1p2vg3BMpIkTEMlHH7On2tJIug/ooDpVKPBWjWO4
Ps7giIy7BoHNeiH2kTPFtlBktqZl6A7jxOikRCEjpm7qlHjdMzHTPWpH3soVIMo14hVatNFZanh6
uTeZHoPv5+fDMN2Ao2KJzpSd/d5xk7u2hmSVo1YsxaF6If/LJiw4E2EGrWuRvrrA94LfOqx8h2NT
94MbS+g3qsrKvLUJ5ZVk7bf92a7MfvuRx2O/EoJTEYLBdk39izOYRHb0gBGxSNTHH34Pef4RcMlC
6tPBOlzs7162ZnBzKxp1zSPkuCmXnC1/8CyKfhq1T+EGfANVUoUrrE2MKjQ4QqE410h6mPTO5Fq5
8SRPMBSQYJjolo0/uwOywo5REQB/nQV9oAldhlIH/o2iONIMzPgriQKbXYWIGkiiAYgCpMl/eAhS
hxU1MhQw5bkR4TuN4erkSJaCe4mmv9DFpTKEjPDy2vVZoQdIt7seAVLLFpBs839VYKXiekvNq6dB
17fZIV/w7/uXcbtJw9On6CUBZgNcQ7OHmaVgxF3GPBcTPFmIiY9owpA6XBgRe3QJAwlwx7k+nwY0
BX1f/yLG4U9Mav0Sfz8f5cepJDLJMEynGCql+O27R7XEth4HPu2CthYGj/Dz+5rCq4/Xo+UEf7iA
DhV4vBwzUszTwl23p+910itjwsiqd1lTBZnXSxPDrQWRS1BDTgsxqJT1z+h/YxJKNzmTCkN5mysZ
mtksXZuZ4sTRx7ltbiHfc5HDracL3UyJ8kWbyrfuz4i3C7wz4AUT1UvMRwDrMaTOqD9CzmRFKkF7
rooJ5ZIFPjwsbVr2l9jTIv6HlE9v92fIXfeuQpfDucWFy1bDlEbX73EUkl5TBmI7NBAKi8BIdnNT
FKSsTNmneoF/K2TxPHVqyIixSSpFW+s8m6dyBYXbnF8csdlUxXroQwRh/5isoB8I4nqEleBp/GJK
uqUBlCtjANA4sadANkB0jbn9cd4QB6kZhilWnJFS86oA7gosH7HuivMtSU8+pjcArk0suXVxlb2I
8dMgiooYvyGHrBRhS1yIAWY/pluQTJvpYPz0xLBs3UOa/QGvmYH/VBnVYeSMzPTKx0EfHhruDdt5
n3OqOC7CUN52s6AkTJQOUVSDYmXmS69ulCGHkMCZttcDUfM5MhhJVoDCfj2jrrJzyzxKgFdbIiHn
YwSVMfmHmBXFelY3rDxL5XZ0uSMvE7tluWm8fAhIkjpCpCEgMkP1ygkocoO9aWpE82fXEkYQJ6mk
EV2f/tlIb1RAwMKiRbZ5RuG4OF9h/soM4eyVHAsnfOcx2GKKFqva9qijFnM0gMnrIH/J8PrcbHFu
TOZ0WoIVH9BccB8vj99Uwn7oznIovkLxXcz9d8aLNhob2fV8nHxq1NAAQsO/Rx7jfOZrMpu8ucy7
+tCJfJnHAmcomWyLnt3St8hi16KbCDYA1r3PGpooAHm+dy9mELbtpfhI7ouDZ7SoScbut4yXEJZk
OpYKH1EFC4eN4fMd3wXpQhb4MSgpuTmCR1pSX+11e0ualDICA3tfbI0lH3jC+onNm3JxtR4hPgC5
AKKz8d01pWZMhr7hr2otp/xcIVHYbg1S7iTU4bYwMnuAGLCz6RqyWlcGDOclw3AYRaNgNulFQ/dU
bhuOXPUTpbxGfmvKDHhYge+DOSFUeY24OYA5tQHXl+hobm0IBZjsLuDm7gUAyDuw5l+h0hVXwBro
/WN7qhJdqA4Q7kwTO3xPjEUR+Zs12vw/11CHq9oMhivAGuGQnZq/rCGnc3S1wFfQQEBW2ipVbkvz
CHgw2LpOgAIqV2M8rZ5Re94zwZrvsuLvMw17Rc2AVarkFJ3PCEWHlIo5+ZeJMCKAE61YAbLubZn+
8DxSnoMgsXKEuBXRnRxPv3vUor5QGRFFoNYwxsbR16Ikm/zxPOckpPuc+l+ZLVKZ+EnhuqDKSemX
e+YEjAilUhg3wLVpS7sYKMIwIkr/s8oY+SssGJMGL4bwCYVqM/sQt0qtvC+b+Y9nFz2IvUvSJsPG
wbBRBpgKwduV0OPqhbC/uRHSTSFKo5tBKVsrNkBOSzfcTNxYDb7jxZnMs/zdkvlpttfrc0RITO2E
XMZuFnqQwbuel329GmxVaxZAfj06d6cZuMGmaCOEYaOoGybEB3asPvDgpbhI+TmhE7E/foy354jh
81a145yD68DjGykmAv+Hk8AsM/su+KPb8y1Pj6vdNSPoFIDFVM8/Il6Mx0pBv4VqwzW48E9gYkQe
0ZTZZwMgrfYjCL7TO7cwsGNzupQfKCz3AfMWpLALq4xJBGRQTFcWvBQVfuoSotDWgPq5K4sV1gvj
fU3P4Tls0v8sPd+Qcm4Km9IbR2ZJQbMWsy/+iX/ekW/j+V18+N4OV6oWTQWyv5vxLJWwU31/YcVJ
EfxG+bBenNo4tyDcDVeFIYiy826vgoCQqP15cMLSe5oQUS5lOlKEdTJ6eX6fYWvtFQJTjqsQxMF9
vHCVxOspVEFEe/PV+gQat/LivBaL2++lywsmd9tUNLDySvGD0CWvaOgZpl2mybjicYtAw02wp9qJ
6RgMhV2PpAo7VTaVAwf/6gYg1P0pLI71evGHXX2GaJeP6Jqc9P0Hy7q+qvX0gytve0s1ITEILqu9
kC+McgSFeniBJPgvQomo2nEmbiuvUsv2Kap9NWO4Fn8GvopfAw3JAexMlGdRgZ5hG+GmsOCPIVbu
c4piQdr9M4ZqPpiO2nlfPo7Fp673EhI7tuJIxugCGVNKG26XQopH67YkIkYNeWNVnCsLqg+JzERq
70+6v8HSUTlHMnDdCWkYA8N3v0WhJraU9OibK4GWG13thGtNHbAjf9uw3oJvap9Ijs9dBUOpfmbj
CO4+b7gWItzAv6AlQEE6FX9h9WBV9rICC/TtBopAArUTNtFMLfhxwWmzKb16fbZgprJZuuJpDoml
DqpXsp8Md8NTgr/Q6N7zusw8Ro0eZfIJv8TDh/ty67XV7QKPqJ0L6Sp+nRSdF7nPBzWh/bT1ByoS
R5Tonez/YDXyOzJhjp3jcrjVMkPyycTOZrwJWNlsMX9IYim5cCdMFiXvSqzzTr9ps1GnwbmDBkRw
WdnIbjLZydjIoo3DaN+LJ79hECcD5lYUpGjq4lePYzwFgXQ9hudMPnq4CeY5d0VYNm4TSJ6QgLgU
KsGRGwzkzPFjNN468ZivWtW5C7qK6BgXft7CwsvSp18jJ8bqt6Edx7gul1subcwKKWkI/ZrcKY4w
B+DbQtVjdVpYTy7I19n22vR6qDsKyoRrVVGnzCAt2OdKsfMxqnicEx+ykHXmMjj/XrPlPWKSiDwx
+nJ5X9RBeLCEuTZeWLL06vTq46RFAaJ7y9frofiaXK1lnVrvdQiaJuoWu+af84w3pQYZEDMl0QFk
3B0P6JL6BmUQzexe8mmnKchYZiK4lDPZDn1lNd8SoPMgCMpoFEwQwoCTO7Qe0x7RP2+qgRSBAwBn
YzogAgRwp4sO45vIqJ9wNgC4MEHou+TN/UQSXKSDV67zoHhUxE3/S1nrnc2uuK2pqQ6syQja4bVB
iJl71YvFawV0Y31pH7pvYyRd9Mq/KmlqkQDyo/wraLUzNO0fhu4+Xj7xmzRFYVEjcCEjZvYGPX+b
/FT0lIBWrPNQm8eClNmt0pmcLuh2qNgm59+znffiCUs+aPaN/K71QgV2f65CcXnebrX2KI4G2iCu
OKHcIx2MSFXDai8GSo0iKB6E5ZwxtMMJO3atxsC5ZOVeePw+9W74AUDXyV4OmxmvILWaFjF332pR
HaFnoHgVZSl/X3N0qxognykQjSmx5EmbmvZxiNOvbbZFzCoIqhn28tt1YjwEn+mReSzjl3/B192e
o4VmEl0p6Grw/M0hkbShdghWlInIq0a++SUP050JP1+9sWWKjcJk9DIPHi4rb3d+PvxLhCEwJswv
w7UiOrCLdpTyQRUjlrfy53slUjuDVJT+rdsoYYBu/GKisX866VsrdRyOhhwjiaHGMepHAMaoKjaU
9EpsZraGbLH07/MV1dILcoK2TuVSW77tto8UKxlYKmRhKbVOoluMLKQv9CrDmHORU55oC6fBlwit
c7yEpLhu5y7wkqS+Dgp9/Sc/PyL4aaeE6NzgZulFBuq2h5rjACY9FbFNzk3depR6Nf3BbYTJfxxs
/cu1ZAzYJIUdIIzOf1wB3NF3GdE+3w3796pyxA12Phbvp+UWjQO3nXGXu7rERBj5rX1pDTFno1EN
8LXajDCl/cmAIBCo0ozmwjDTsLR/Q21hu6hjapkc+RGsfsNlKYspOL3A8uOdueVjA9Oru5iW1fsZ
1bbMKiHmvyNCqKL4WMgoZSlmpJbBn2tRbrsfXPhORm+jzf4hi7JZ+er+npR0nhARzYta6H0SRNWO
x/5Ot3j8vhruKLk+v+z1O4f/H5lM92gnpNW/Rnso7woxM9FAJd2or2cAYlXnaPZeODz1rGyhj4Ru
QBmVEebeZNzXlkTAuvJjp9yUD/DuU0g+5RtCE8nwcyXp3Z+qLwOoD26+V3/xqLgXNs/uVHGTzmzM
BOyD68xmNaCpsNxJEmnf3sWgJnIWtBUujJIC7G0GmkTXC4RrMQwbGrIWQmr/ZHfC6AAh5wTsVWwW
cG6+ddc9Wrh8rn7MnjkLmT66oLx3apDKCpGW8mMhFAV2/FuR/8p/6VIUiEVtCW2BL0Qblsm10UtU
JSIMjcC5HE7ne9RDtfg1PwUJSPpwM7jIrDorjL6z56FPXCxgl59FqgTc5ADTa61JzHQKC4b8P8jE
X/grGrOeXXDw6dGhi9pXK4pt0OxCjzTyVjqcp/zwCWcZlpJrpJ8tQr49Gk/XEjcVzp7EPkwCmCWc
05kDZD6lrVOaKWqbg7yAJ60FebHjaDOpw5VH13Vy9F9MOHc/cfRbXl2ShdbmAmoThREKwe15FRMk
kD6z0I+OgR+I/Qg/Zh+39Tf92ntybbM1T/6vWsXXDcKPLJLZ/4/EZh0Bbq4+sf39ghhCOmuafehw
6F+kh8RDTkQ/V4uvxoO6UEvxMVsS26tzEmfsoXIimGdln0MQc/18EpQriyP14udmYVm/UpNsQZRZ
x7Aux4ukiOzzmcS17+CulJFvqoFt+c0vbkviVMWGHpD0MXyjfjVpT2R5QKA5Xj3JS6ozep/UUOBp
xyoHQ2u6sYWjLH0ioqdOapvFLKKqn+7R2EJOU5IPrJhoOycE1ZzwU/a5tMC9fFf5oslABREeeftC
uxiu1cFV3piOfNBwzk8taaqdTaqyCbAyarPuxaShjlZcGXo+Geb6a9+173Fv88nDw19Wu4RR4Oxk
aLlKwEzjqmcY9MwgYQUmQlTJXh+U1MfeWmv4TdR7SKIOOL1iCjV+NLGIIWOXbu7GQc4k4B+92m9M
cwVXDIqgjXdRs3V+9j+WQYvqfuuVQZ5tfkjlrKy87F7kXjmR3SbRYRuyLPAgCkDKmX9ttagQqohI
bxIw8kvaWH19keDOOkYedIDn0fg21dTJgPkn0iJNHV63OmSTsmA9sHY3rHapb5Y5q+UlwZF5PY+L
p1eHnR46iH4X5/asp0joJkfHD28fTMhbUThy3QwEb3UcAEUezzV7fLn/mviaGPWJTMOMJWC9pBFk
adhuWSYWfg7qXVC0t6d67RqDaNuINn7GonWIp2p2UvwmFLyCVaca19d8nKsBWKYRxYOOlzLmReTK
G6d6wPhtK/ytxCnaHPDkkP/FxQoT0O4FwIjwszjaXSKPJR4fee0V4Z5k2SMw34x2LN9y0NcFAIBg
baVtVB9P+DOKXJS964PHI6e27Mym+pOqoGThVcle6qzDeL4QmQIRPA8jLp/gwSmJZXINoL26SEYq
X/RpLD8PlpC1Xj2EsL1XCeonTUgfLw9VTtm/5/9AkQOsQueHVgAOlAKl1D2YLUE5FX30rZPS0qqE
FcTfnccFoM4tq6hvFONnqSuQtG82YOwxfKpAbKJgH6zVWIIY0jyIRzQTanto8/P1ACZ2f1cgyzxs
ekcAlLuU4Ql8wHhjTmsLw/71iZYPvgMI4NE/lUFo4WHEZftAKM/FdoPlxNyxdGKl6mGEMsb2SCfl
97IlZu/195CaD0BUqPAVnhd9/9nj7uVfZQ3jxl2QWImB+KJmjk5wWEYOGnP02lO1avfuAlfoCyDi
o+7KQgVuG7uhAWEJOwIb7UPidYJ6BXvtLOyYWkkXGQjMO1VXwxNWJwD2q98+AjKfsIpKZbfNCosy
BZmqcxm1iopbDvEX2Vq5wTQcjAAtmX7PT8TJqJ9ak8wzxSKn70y32cDFb7jFLIvV81pm8cYZGn07
9aPqCpfa+me+eFHEWhrgPTnzI0g0oymDLu40qacZgAD8nJ7ArpCsY84pAqvZwESf4Rf+TJUPedLl
ytEkHtuWFE/1jvK5HAqJvQ6Uq8TdEWsmdb9/zx8Xbk8o9raySlZ1RZapgU+7oMXWyJ/WKENqKGBz
OLmJPa61FrQIywO0c59QX4Sy2wnQA/j11wu5lhaOBNK2BxPmW7JvBS/sGtvTJkYcgQXLhO70tMLl
1jhYz4+fA1fKqUNQS9SxbPFBIiU8N92sOa1LAqVahi84zNbrYdxrSlKcJhdik7F/7dYLpwXh3p84
lyCDO7pIRT6E5O2O//bKrOwvW2fsfcJyjd+pUPHUTDBGF4P4PuHczcd98APkShFo0Bd5fpQWxsQb
+gD6xyURwkzwfxl/R7Zcfug7FDLSSEdgi+cAwKuyNFPEaLeVtVqUtqHdkWi+JYIqIMaPv5r5Jq/D
b91F5T8B5HizNV9l4J19kNZgH8pTUGCshRra+XoaRp7OTd1GVnvMYYU3D6ReoPaJPtlsl+hTbhG5
RGvyReGaHKL0PNweuHrxPG+tCujMgQu646axJ4x9RJCvKUQg3Fbbf/0wA9zc40CX9kVy85tEo9cV
Vt2sGJqEP15VIlbAymUtGweSDrQOwdsPlOuJT9Dh554txjUxk5UlxoTnlugM9y7H2QZOJoVW7VtN
mzo/HEkm2tBG+R1gHGH4QpT0JhVaYWCbEpSzj5FfphtRpXzT1n4tjy3RXkF/3lYAj06vJAWLb+AX
u9rFYUl7wYeHPEoaWf844Legshqj1k/DWBo3JuMrmrXic2PjJE1UnEw2qafbZtgfGOspncsWwLSJ
nj3ut1hZdG+kDYVAicRwKQZ71aszRK1H54ijKlWErHhJv5oJ6toytoxB2vj/5uux+kV0oqaoFKTG
TBBKWkdShFwgGrdCIjdUNjfDAfWoXiH0V7JmxmIMCyYl8gz03Rvgx3uGv8E9C2d6xWotrIv3BQLr
OOJC0Dv3/ei5KcJm3ok25WWX2qm6vHOLUXgUfBwB/8p2cJTr14c+2ISlpxBq2Of+UmmxQHN4DlHE
W06GgJm8frpQpz5emFokvbQwVwJznSeQnzOIPXIpuYY5EcDA/EnORZ+YcRiS8oWs595fFm/x0vlC
RU+G0YHu+qq0Wf2ETCMBBpffD9J7SFXG7sH70sVQ1ZWF7MpdFumqfq64TTDu+DITg04DJe2to7Vq
WUX5y2soLGINaOn967BnYqHmurNrf5GIUwLq1OqWIwvcV+vGumAy78zcOAbkTyTLWzl2WHedg5du
Ybe6lU6cPmbVoz5xcy+MYsfHKXWNJyKmfA8+571M7RPWXHkFalS+uWKsRJ/zwEid021Et0knQ3Kf
S9Edyk2OXmmjgmPk0bW0PQ06OYBeVIIkEmBPNCMnnmjcLA9MhYKa/eR7kVK8u3PHaV4gVw4ApyFe
EYZxHBPrslVbiOnAQL+/UOh9cPn0WOu3aM296Ax7NvGAD+Jijjct/121uRgpOgXnjosM1ztUrOsQ
A2zl33RXukaX9ZKYiYf03mBNz6GXPjU6KnLk0TUvfzmPnbCcU07e0h0l5iBpeVFxYFACIb7Y9iAW
+P3Za/b3ouiXX5EprgOMHxWaIgo1MeOe5fWFO2fyZi/MCg6TdC6v+BDR4XU7ldBGPoUowHtjcoWq
OtY/BlHIh7Y3C/n5Va+M38bkch0QxJErp0y69ty/pXMRNzk+gNZ7CBEtHHatjajJRDiz/twUl+Xa
XZFbk5PRCSXAIeX3QXKBtvZ+9/qMy1QH3Y0ebe3Td5qsi8uX8esc2x28Z30nG1aHD6S4ulFSZT8Y
wBILirOR1bzQk+1h8H7J7RQvSUc/AttI/xl+armSxWLRSU4vXQA72fTyYtZlPRdmGWNobpo4ccOJ
q/2eXMQtDvYRl6JRKF7cNs7MXWbGjWm0h8EPjk7CLrIsNZEjc7GmX/xSMr8si2VPJkgKJJUrzxci
NowRIP7nTMoclB5r/mb5c596Ws5E6XG/nySsgY0XcfCklOyCEWSyZhteNEm9DbJ3PVdtsJ9N7dZu
/HzCG1hjmZLWX89mm+A1sjjwiJvy8ZarB+/2gpW/tupkByd9mSqg7bWSxU4dIvm6oP9ZoV08tTJ6
I/w26hr+n28AhAHKICNZdyKkpJzImzuB84bOT29KoRv1sChzlnHxbpd19udppRGuDRUwHiJFOEJF
LNf69yC+6EUHdhtM8cMIxeyqoTolz2hdBNhj8l46+WRaGiVcBnpcm+0OUbT6EkmQsiYC9yEDYl/Y
qsssEkr742hW9zanB5CaKfmH7Ekajv9Sx05EGNd4hTIzqQoEDJYeW4e+GhXK3WSNXwL9ZWJlmpFC
n0NMSRIpU8rsf+bsrIVRcQzrp015XQ9woziAAgIO43RO8sbcB7nn4Q1BQf38HWP9GE/Dve+xEn/x
5gl7e4lt6+WHDKl/cLKiY45AMGruiADastVyCR+fzTMaK1xzVG3gwaWFA8IHOmqG6ZmK+iCHr2Gz
QSHiPRsAyMgtnmA5kmK0urXJUjh98MwiClWekvi1At/AdVE5HBAUv10I+FLy0a28I5D9KxvIxaAi
AvSPLb9HqfCNYrumq38FKOBLdmmCUzVK+9B+ka6qxTgHttrJx0KGt4w0u3xBtqYF0z3UEzvlB/Tx
5AEj09GS4CCQrC2ADCD5agh9weWPg+yruNbp0RS+pN0BvQj8Zb/Ldn57xN+fjmJXwECGbLMombOR
1WQR4HiyEFWgbekxhv6XOc3FP8Dst+4cUEb/OgkDLBLIXh/UWKZGmS9/ZilVrOMT+hlxQKC/b2/4
k/jE6gUQtxIeZuseDUg9q1Pe1aGxYNIKewmB80ZPcDENfF7tx1yQ2Vu/dqXZ6xLUH9mz8/4n+0cY
Oyx/6DImL/w3Ha4G0bB7w/HDP64ZeiS13BKVkE+6oIQWQov/Vb1hMeiBvRw85TnV8nikBmqo0vDb
+HfkbSjPw4q7Ucmoq4j4R051Jvz6IUl0hqPD0786x54bYlhCD9ggxjlzP5sksxT80iTMms6Hdm7D
D7oMjEhHyhPUSLNU44DfhHW1QP3OrjCgRyI7a14RTccQaWRia8meeqm8ezJdMnMLUUpW/YGonRVp
ezJdfGQ8rDcR/J0tl391But6b8t37PSEJdZ4T2LNAgbBh52hnYGwy6HfgkNHKw5ux0q5Xi/sub00
MIvM4h7c0GXjc++hkzoHYPjjlErnXRx26kLuX+1Jhj99XpRZdxYuYJWkxJKx/Bk0ltmgbTqDJS49
OiF5LYVOBFcXkWtbhU5ObZashbshbr397+V86s25aaGBckY+pKJDaUdlA5pPXhm5CpNG6Z+aDyKW
wiQyI7D/N73TnzuXvbsz8NZEreywtGFoKOHb6Fvlg+ZsNk48mzTm3U4ruv1AJ1jWIc2DYPtss7PO
Yi55TQzitwu5X9CKko8+Eb13BKP5ySHzhY0D6Qg2UgKOd+HIzVhz1OI9cSFonlodoNgJo6SKcEoY
OpL0yzK8mIPoBsJMXDDGWmoeo3c6AfngQUvx3ZQsk3d1y49JjdpEA2oA8sju+pNYWqRRvieBO+O5
UAUZcXf5xKbCc/WW/hlcgsJz0YaUMmGI8vCcY/DDJ/GkLOmRrF0ldwti471gAIYayiInpV5RN6Hi
K5bC731HlHEdMMP2rTRq48OARqriT4wjfshiE9DFxTnWQ1ceKmIXN9dlUn2SLFJVdaQ8ETZ4+Svz
oMiawEVqyRBdpBNbk5zZakF/XuDAKRdyD5+jR0rhfNZ+aZoM6bXhKmuGVboSXg2geEl845JIT6Rj
gG9HqSr3iGi34YAV1hd1yRNG2Wm0VljKjN795Ps9gc+A2pQ155J7oSCAqoTwiT02uiCgHgeqcrp0
dDu92GC2F8+I3uX4tFqbdOlQ5SClZXiARe1fXg9452cCsdkMXfuA7Jv3FZpk9pAF9vGutOdlhaKW
gYaIbH6o4o8oz8/eLFH0Jn/KgL9SfV0fQyGJvtw4pWAy4PJ53+LP7W1qG6Hc0g/e/JXxDhwZ5MDY
iplSCuqdK5ct/rFSrIEIwHyVLqoJ/aHxf4n8O8vwrhQPFiVVBKCV0+ESgeTmXW/gN/ZoZgQHet9s
7ClPY2HaeFaLM3bIVVceyiv901Y9Dum5x8BMlMQAi9d+ozKiE2kuVo4f1+c9wvmIvFxF2mROz4In
jKIt1Kdoft0w/pEV2GPwMIERtFuYLucFAudDvOQQp3v4fXNAdtNxTqBN6GG5JmnM9ivVAoHIx4Jn
VVzQ/Yi6YXahZWHoeF9LkodC8eYxt5J+T7xnjgojk7S4hxYlQ8dVoWuW5cvmIF1p3KP6wS3wtDCE
qBY64qCGwtzXv2uobwcK7R5RSuhsfWSuS8RIx1JxJNrecEF+o6HO0bELK9QHsGj/Y1o6/O9wLP44
gU4TqU9x/YOIet+pkxZneZquwvygj1eimFddJA1rjwkI5EWWizTj3peltYd4e6RETwQk2SghPqoz
zrycxKgIEUFHPoJjLwIQaAKOdQPC5pxoe0RKPiQ6hSzV/Rj2Rlv5c+xdIc0O2RbpJZE15/StRBb7
ocdnV44eQzSFuegfb3xMEITtctianPFxf9xe31kZ4hJEGeo9hDUuopcXT6NpexvIBagGTkqMZA1m
McR2Zmto8urlA5pMU2uvUAS3sXUYoUzUW70jfPiEtRRTFToO6bewWUb9cSLcMRQATDEdFSg83P7n
4rNzpb6ng86ATLPAJFzS11FB1lwhh0uQtdhQ7qKJSja7Fzm35FVD7ZqgMUasW8Zibdty3UTXDA+M
fMos7Fjzi+LllvzhPI6V8GId373sLAJpvWnkB+zBsYlKkBbFuAgjNptKtdO4aAvepsEn7qT7s7K7
faNVWDlDouPCkpOMoAYELHJGeTmHlQfv+U90C2m/ghTo8lBsIYr/+YfJdO/JRYHPOL1vakO+B8K0
+oojjkzoPyK059yO3E/BzlmDY6QTCDHCvtT6lxccku348Q74+fgcVfg1ou6LOfJIYB3bbHahjug7
KZCbjx8iLrwdA+gz5Dz7EYw1Sceh4g8HPvdvzr/jLYF41h0rn3iHZYCgI/v+ak5/gE3TpVVLObHW
WyPganorJamczAQCZg0Ldcpyxush+Xxq7jY8YEBNb6nmjJtPHio467j8oFEor4Xmou/sykqxEkbN
bor25Cp0WGZpOX9Pr0vYUj+YjQsuDnkpimxlzbqPpt8QrXtC6S6nxrSgrg2xyJCPfymlviDMrS/a
/2GflPM2wyKghG09Xcox3M1OR4Sn/p3CYvKg1DH8xOlMog2txFh5ZIgCQ0P3sS7mLJ2X+cPJ4bwa
2Cnzy3zYowfkaGaDru5NnmPzPZ/QGLBH8JBRj+znrUbO8L+YvSMa4N7WyPy6NGpKFpDTXIIxhBm+
TVu1xqSm2Y9wU8kYa6WeYJPS4Q/JXnYcypj9AUxAQwprQLfCzOp3LIh/Y64NZ4bxy8Pc+3LGpCYX
QoShBTbhfhki6+WFhzc9NqH5lk0cUK6IF1xYYrIhZrDDZWIYSKtd21fNHZgeUo5PQJ8ltKSelAya
CzoWyP7vTQrN89wWk4Esuh7B+o0Cr5A3qbwc8I6u0C6GO+2Y03xpUl6dmFtl8IGNOgfry4SgVYwh
Wiq9QC6+NEq9/A5xrDbN5vKLQrl0M9bdH4JhL+yEHJn1hvyWci8mpcnCfXQfiO9edlrVT3CoQ4FJ
uFSFspErMUKZdFVZ6mYpMhJgF2B8PPB70VFOwyp7PeRBbE6L4Np8Q9c+d1jkKZamOQ47kxbESttR
PNBcvaa+AtbGXEanVEYpzaWKkwAGpwM7TxHRkZtqlBJZkfjege9/CXs2ZB5vlrmfCr1JsDmFXvoc
CaKivcgcvIcpfXGBEyFk846LdfSLRehPn8VarEr7mBjdytXQ5rWa121kuV0jj9BAgMd/n9KXt9CX
FqaJC3lv2Jbq7e+xv6yhnFs2kVxqnMG3MNyN8nuBdewl9oZVy39FntWD+G3z3RR84yfHXkF4zjwj
wCx2kzg5gBMianGg9kWYFhxVEh3aPNPsfZTUHmXMAIYGWMHcGoav2GPSHCvnfer4ImHJu7CHDuBd
PkkSAmSOOvDmPkonBPbsz+N+q6RULFckRzgVlXejjKu7NVxXOmVdm3amg6bY/ik8+HOsbqIsLxzE
LX5B1Ivp8XGz7VC9SYFhHfAX06eZYg5Flq29UkHq+ddYeROHT2uBX9Q6zhZgYJyBzzxaxdqRCvS/
W4XuN6kqgXwoiA6JxYC/OQ1xL6JLYeZJpc1VHKVA+1h5keMd5WTYUh4qCv4nlbIriIkL9FXgfyqA
S9TsLo1ZEqZgVWvTzOWIDz7KgrRf53tF5nT4UHJiGGBQT2mmeXeR4cpgtmpGWtp7QGbpMYxU1SP4
2XXJJFvKtEVUpt2chWNW7j8S2yVlYGIPiZ8b+z+3xcInndQzBy+2157Q54n1p0ZgcGZnZdFLQfiQ
qrBt/j2iAhdznYHTG9BKk8ad2tp1nnIq0WDPKuzp6tN8s4x/efm0jIkhBvmKnPWN6DRx5rWgnhtA
iS08eBIGipwTMpQaOABcYIQdPvTUUjS/g9vMAX1+aqP7uNUIYnGHdeVK37hPDtuhDzzR5Vh52gET
mNyZi7d/cahmfwVxWL+ar+gR6uXUMkv2toUQpKHt+4RH2KU/7Mq6R6N9OHHyarx5do1PnHdskxPF
XuhRp1OKFg0kN/27qB64u0Kur2ZJzTZ7g6yEahObZPH3sBbVQ4Mm9Y7H34P5XoeddAX+I2X+Aa3+
hkROFe1rQx6x/SPMhU6pe2S9QL7t9rm9uAUbej+cOGtgadRVB9VKurgfvPcvDqgAwP7y14mA3TwB
RLm5olRtLc03a7lixp+1zIYewdQCgdtytm2aMF+K2Xfl58ii5IfZn1oU+Q8I/zbGdappxG7SwknK
dENVA6EHlJsT4DKsGusvqT9+ohukg8Zf2EIapMC6bHxKOBrlTHj/rcBbedywzp8pLHgzeFunwNg4
Czr62sKlIgC5EUnv7h8ljiLLjYrwczZoIxwLFp/LIDlQPXr3v7lK3IlrDqj+pgnlbe7rtvnudYTk
NZlR8B1mRyr6P62/ibczfRaj7trDgco1pmNIyfNvg/X3Q/nlcaHlWi6CS3u0GEyb8ZEEVjALHR1r
umG41uIbLMJq6WGwfy8GjIgHsuz0M21sw9kvN1fhtV5uFr4YKJhT2X0Li510BBoF2Y3S3y12Kn/6
1sID8N3h6Es/Zasa8EsPpQySwgoaB8GSNsCioQZyLwehpHctweh6+PFIMSIT1D/GL/VyuCo/49uH
Sw83erLPaQ0+zS9ml4bAoTUeEIhryixKWxVbaanHzBiD98gRJlODevReVBxNvVFMTBhRIP0avyGP
hSU9VhZVHvHnFs6R2nbbeDxF/gbatwe2ciuxOLFdp07VM71fnzINgNfVfLMtRGW9J05NMTeMdrg+
K76esbDI+EmDGxZaEIubp58IQNkWrK8PJHrEi2+D3u4N7aiz3HD3yYg7WIlHjLoKpk6ON0e1qpds
LfPHxlt39CsNYIX0DGL8i0RHK+bPD8Mo0Wr/b7yA/4lrninjV8Xr95wYaL+7eu3gixqadgqcQzpo
wSPTznIBgVTlnY0VMkzBeCfQILBsPvggjfLa8mttCu0D1fkQT1Wi6jjTHT+YewQfMgRWKxmvcC1K
yLQb1ww1ovn2B+lqQY37NVr1Y85j8AauCS76hfqGeN/v9eNY3Jb2t2hvRMBGQiHcFnsmg8tqB23/
NcGb0nJQjUt7yhAZwjLLUGFEYjOO71iVJjlKns21gZ4vv2CE7EJzPKtTPYT772ZZpR4qqmkvIdwZ
Q/5jQF8o3gKexhZcl9wYpVwQJLUYn7BatYXkc7ZfR9o414r5P6nocgWQHcK7MDryNRUo7CM1MRLc
Bp6wyy90Wah8H3HXWNwu8ATW7Kyu2y9qMefdM9EDlZvFvkpzxiO6rJtdTJuacRN7hc+jIVDgY+PJ
alIEhpW3r5dxhce5qHuLgxlbr2rcg4Ka4BeoOSSDnz29TCbW2PcJzHPwk+0jcoFrv18ZVPMjM9ip
CCHNkFvJ90zQPt53pUJV3QV4HIKl+mwnBaIApm59oXul8bHGNmPME6SelrEwfLgEbbzbz6pa9viv
mewS5oJiGdCl9ku10s9f2a9o2JSnOuO6i53uPH67R9f8v1tQcZLy6SWSltE5KElOeyDSUlww19sZ
bg80/8/ADNnwHi3p0qebHINPQFe1DbWOgoc4ruGO9plohZ2X4VHYm+SQsdfI6liZnElTddH9mVRq
uV1huPeK/Ig2Vglh2P2XyOFG7kOMBQXXYKJP6q3Ah0aRqUKXdo9Zfr/x7CebYYYJyL688qs2oVIt
0kHv4Fw/AqS0ts2MN1NsqYV7b/4fU4b7oZdCVz4k/QTLCgNQsGv+fnyVhrV4JVaVVOvzdHZLlQOh
M4e7xJgqoi4xD6eEl4HrAe80iTydIHmbq9OYWktqYPWjg6SS0b4oGXcDI30hQVnLH7pm6hdbLVo8
b/76zO6Eaxey8E431OAVYR4MkbpV0Unr+opZQLvv21TD3bwuA/9FuVJN7EcPhyuKlM0crShMEyvE
y1gGm98d6GV4NZsDySBSvxy7XmVsbf8/jC5Z4fEM6jwsE8Dbfl9SvKpaviC0fgA13OEpdbqtJiQz
UdbGe46jJjy7Syw4YMoFbZvxH/LDRSKzlo8H6ZIU3N1JzTq/X4Iw0CNKxE8p44S3WboNcD/EFWoc
PwiHoi7GWQEy7/DtNXjy+8nR3tT9yHOO2jBENw3qixMvf4sSAzRivuqpdlWvwKq2SPxeY8xPx0HS
W30Hkx14kxvs8bySRnZZMh/ZZ0s0caZtDsxfz8M/cx5Rbw4begZr2lgpdpV8mLZw34trZMkkASDF
CxBxny+uGetm4o0wYXzTcAcu0Q50CQRSC1bJHxo7oe+Sh5GV7weTNS6bzG2528jttFp++pGwtXa4
CXM9lHFU4WmMpACbT7z9x9eZfS+rBScWwmR8UZADfLc52qtNZ6iXdWV8ygVwl9fKdbEe24RLWuI7
CN1LAqynY4skhDaGu5MP2WRLX+kOOSENSDbHO6tZfAe68Tz87HwnBPH50EvHaDAA3aKeLhmz64Qi
PYd9R99+IYy4dBv1HqJzHIbyiZRMYiA8EnEyHCB0/DiSaEyx71dLN6uVAYv3Xx+S9cWb0Dv7EWgR
a9tsAFqTtUcgAHIFTEJ61gIdCxwOvMyR5rEz8lWLhQWgaoB9BZOAwF9Iz1vSdqVyHDNhYbFojkH8
/5Le8Y01uQ+pzofYxRW6TUN19EnbQK2BJv9YjLRIF5CUojfBgNgwQ+td1qwDf+wrJuMFbxznS6eJ
f8/qvY2BKBs3SMlb3ofquWvtU9/Xy/6GGrE+z3LN/rItIjneLe0y//DvD6tTZrXkZyemR79/Tg2N
eMnt2d4tMcXYSU5mw7zdNajZB24TdIWp88Eqamlk+QJBdiLOTurMCQe9lx9tG5XDMSNuKQpR9aot
eVrNwQORm/TZXJ48qqvYOcsbrSQ8AbW4o1mXcqnUMEFCE7Lpyx59rGeqUoncIKmfACiGxartXZpL
hPSI54Ca2E/puqe9g23FdGSQ8gYE+HukUmZeqY4s6AManiT2uhbOdzUGzfH4Uco7t0HQbM7vyyxd
RzKjzXR69lhcH0iMAsIg7m7NU6ovscgac+BCqtHP22kIXUQ6hz6qLRjoBLmRj/bo3UQGu2CRUbOg
qBNRN5hekbyhSolJJo8+5zYe2Qeh/zjpaXonnQWtdKRoMyJBmgbguZWHtzfnqHwq1LG37/mwtiDN
+DR8YfdiANAaippHdnPGKKrq58mB1P+hrKVVzbrJ+4WhuN4LZGKPbCBDr+W3COODRt+3u+IsdnV4
VS6be17PNfCA1LujVkdvFse7bcb8QvIjaZ5Lo4KfUxlBC+0+OzK1KKgJ0yE/xZpq8LcTqv3Vfx+i
RZms5J3PTvByFs4qsKiNoWDSisgGOquPcOt+D76Kn8IXdqCa1Dg4d65tnbRXmLrovuYtIs8ZngDg
tgpf7dTQjhqk60tBlJgTbrQe8ujWYOVx3A8BSw6idQKoUshnrfscczaH9MtVVjYC4p1mj82VyZRo
NLLDQTU1rq0fvkXvs3OkDlig8kGwBz58Kj/hSUkw8lelcSwqh8m03Jxp+Myv3MD4r6Sna/F6rPim
5rijQnJVHzhd1pyC1vE7hc6XjKAtol9CNoeuTfQ/FEDhRLQSz5TKKNcuf337Ora61t+Ph4TNDpyQ
9ng4GH9yIimaBEPLNoe/aLehYEwfv493Wc9xeUI/31ye6n3zML2B9hsz4bmsL1v08fl61tv8f8Qj
eUqrTf+y01dGb+2DiPknEe0l8EZdoujfn/N53mpcQA4s1hpi5nmqNpTLj9QZKVMu2l6FvxkcYIBv
utN6LJ1x7xfhe0wppvL/u5aQme15N8CZ4yoJvO21CmGsQIS5eHXvKcQyZJHMrmqb8CSZcvWqwNay
4xvjy9/fH1boablH772oCqMbLgaYsNl4t41F2e99rrvXlpnF6st9fRpFm0uq8Q7F1ONkJdybHTWZ
1iB39kj9NNvYESNVAMFdYy4Tzg7l89Rvoj1deDcstNgWRSZACNwrDHyYNVBGk2VEj6xFcydxefTa
7W0DDwME5WrUfy6/O1W7bztK/NiHoZuckAmFIPSBArmYx73fvHgHBGn58A2salYAzYcIMHkR88Tq
V+dA/PI/dh2YL1FPPovLEX1p+9XkkElsLwDf2i98vbPAtJdPKEpbnVLmiFDyCIaq08pfg5mA2GXf
I6YdwUyGFADkznKEe5h7EOiTW/Mm7QvOIYzmEShcTa9w7W420o2MhgICP6OCbUOmDCy5+0pQYACE
67CwBMpWNTUSFCjBcBHS3LaO4niDLrEWTVrtnMjaaSFSLd5GOZlktXYSts2AlYAWJqLfLRqGJQXL
P+Nbnl3s/5JXrPym/x+fLy+oNxf7I6LIL7EbVVDs4j20o4Z1aFN8TKOpcPa5xK5fGwzYj/RNbIlS
2XVkDhqYk6WbkRSZ08sELJGedtyJjUMpOO7QDLv5Bz/nqbm4Rcfq2pDqVlEOCjbAM5NG6oz2ah7H
WRSkHOcFsCKQiKf5Ub2wocYHJZYQ2seV6Ux4iQxxP0UkjutwpDJT5Hhqm3XR9NtzE/mF/CjYKS/N
BaHPK4CGOcmu6XPf2owhVWTYgX5PGdCX+MvS4fSlpPk3ozqwk/tSiutDmNRnDq4MawQHZ8v45YF4
RQotJmXkPjsHRoe+aHphQDDbaWOpEy0ay9fgrAD1dklun9cplERkuehw9t/J91PCR98jxfx0MTFG
Q6DKDjBlr4eApC/hpdcltp/uVMeAp7d9MShdI26MivI1a0PnKHjmdfcCb4D0AIxofpjLwXhjMJ4S
gRiJ47fSOlHALUWvTKAb+2FQyY9A7gkHigCshKvCdgPg+FFpkx7DLKlgBXZBBYBqu4WvHxarXew1
2rd8ECuQOm9V5YKyeo2+Iu1Aspb9SlZ0YbUZcBB+uzKnU2a03AIuGUAGoR4/PPLrqEKi1u2Y4HWE
HWwZFgFeIuQO4UTibLg2XhaXau8OnhqsjIDgHPQ00QINRKWzcppkRx0VACQXowDYNXOCaG/ZHoJ/
xUXCBGYsR15yIYiXZ5kSrc9fQjh2SqvHjD9/g1jFPRJDRukPM4io+Erj8w54/sdHmuECMcc8MuI6
GLq56YAIFBuflSv5k94CpHlGuQ6VK6oCw7V0JoAQS9S88Dd+l0HmMez430qzwCPyPDnAt+6nTD77
N9xkgAnzq+bfG6nj82ZHUxCZrBUvwXghDJzXHWF8oVXj4wD87sZBGO0NUUuGTulBbb/qxOVX9fFt
hrL4qU7+L17dwc1v2A5n47o9byUV2r3FFOzQ216Y1Qc8AhbtJM5x8JNXjB3YDetFVsHL/k0HT9kq
V4UnmLj6YNL+DHTVq0KUxb5F+nKw1B6Dcc3dsgJAjgATmTPZ6e2L+tssyCjehsxrbr1D11cYenku
ORhGXZfbPcBpPczkGkZDUKyzXeGGQe7PRySx9nOUuSWeJjI+EVlKIxNhdIKuOrTwRe4z4r4g6Asm
VYbjeGZY3+YPaHtLMWXKlSl+x8RDYUx3PfgvBFTKduhrrnmmvdRAamCcU3Ov+31I0tIEp8OK7zDB
lf56olHpVMnmnzDYHdtO8d3TCS8Z7bfICnv03sUhnINf3LxSnPGC+95tDFaD+oIEKPAOlb2nA1D7
sOCl8KHRWVWWut55dvgQ3s0W9xm0pNBB0k5NHFQUxVK5w1GbcyJJGXfLXDTILr0SgP45mbZxdr9q
sbfvUVd+zc1FQT2lhO7Qu/gPLlGQ9drx9ykvOzymno9VGVO2nehPwQph0dAKwXnE/c+xjETuOcmO
NsxoTipXDta5Xk+D5B4WJ1Nblw9hf++TIbHjhlhk5iQILc6yMLsSTOGW04+DnAdG9Mk77Ozs9yVZ
dt9LX85xx8IL8N63GVx2XLLai2dUZkFowgmtdh4SALNEZH2W/Nq0nOCN6ltu0aI4axS+X6w0aUa7
ZgLpDOo3rA/kifSAgVi4Hy8hJo3tX6PrukdVkh0NE2SE+GTQj7Z419om9r5iR66hnAeBC6FQeFEG
MCrSVTt51/onh9gSzd+Xg36w9GqvccIfNM6G7+bMPmzN965J8VrT61YKb+QLDdzJc9OU0PNpAmkh
Hi6YEaSY8LG9FPiU+XTUaw/gP3OqloCPLlAgv4nbDJsLhn/+6VZRUJ7AD+RCWdNdxB8ZQ+pQIkwV
Mi5wHTnn7XlZNyYWVHxNONMwRGADHdaXWi09Ha/rZ1CFhM4nmeDazHUygSLrM21W7CGKleZkOMKp
WJkcB81BaobgTYNqVpl9Yg18yzxLPuhX3tTj4pCAfZF0HKr4JkS33RzbGzfavfMQQnRjpfX9QBEH
ZV/qlBD9qNEwtBvL9/PQjhTtJTiVDDi2WYldf73XzWdO0RaOtZrJw6WYPhNNhvZlntgezEuV+AZ6
sim0fXWt7q9sEjQILWskJxIBoUPrdNKA/AyUIOSf1oQRPy9361xP0oE3maiptFFGPxWoTmNd5RkR
pDhASXP5nX3U4yUua7rer1YEulgUAUZaBnoZ+icB/NPf2iYOJgiSocWx2bzWdnZyOETG2VyJZIYJ
+W3g0SEuXEXXCw0CZ5cdRH0wTyKHyPzdBh2XFW+YsGUtG/4aCo6fpLMA0H7mcigLZtaEkgFxFs6x
k8r+olY59cUSQMReZhMkge7czN9S3S6+uOZgmK15MVQNNGSc7drDu7eHCFesMER28CfXwLaUrYoR
G87fM0A0Q8gucJn8nY0ARc61/dlHnAbe81ePdaVrtdl/gabzuSJWaiUpAqAS1nLfUAhWFw2DDTyl
9XuHhfxg5uICMwFJ8gTccXhZ/mklhPDKg92QcpwQyY2S5pYj7jyAoKKzoxO1+mjyq9XzXUUGXMi/
xri+zU+rl3NlxPh2kq8CCNZvwZctGPO/9uTtMHdj0SkLS2oyAy3+Esn2OiXzXmvikDusE1iXQdv4
EVPatNQBdCXhwDjy2RLdhlOEZ6va3pm3rC2GsvEw0XTiAgABVFXImFU1HRN119Wi2DvvJ72S8o9l
5xHpNC4tVuNyS8TBAw2MBDB2v8ui4mqeIBI38anex2LnyCyk8MCkGVQ4GyOJIRmbI++bhmDsKkxM
M59vacSmDpjJ8Ql6JBfjrhkFynGZBMUvQ1nafyb5T8n1JBtIn+ob22fw6z/gxAW8OZTOVNuEYGxR
khoKdGzzBUq6y13fU1g14vtd2HNXx0zR8/98OfF/yvO+WXkk8pzKz+7nNAoefGzM54plaaei1drN
uPBVoiemeDe6VQUZdxUG+DgorcPulNAWp4PRhZY5WtyxXTYIE1BZfk+Lx/qTgePf2Jp7da78Sb72
HxZUk7DkvTbkdXfe+UMZAUJI6gcFY87HCLg5213Q17yKIQs0tBdvBIQr/HaUdKn8zEdmmUrHyCx8
VSXH5w073Ke5DAwPGoLc6khRgMDts0kMNj0uYnSK9SQmG8xUC0SPJWpCBYACdkxqR/ZxnRyzlwoo
YqOYX65u006/t/y9XnuTqpAsQGZOMvV75FKpYRqjn0ZkqJ+cD56V+vRLvGrO+1ij3y8MNKCgbNFw
SbOcOgd8fk3Xd4CeIijXJkmqTdDTpZCaXOvkbyq9sNhJ2VfO0uPK4rxW8IJipUkaErHs7kOBtkeQ
6DbHizKHQvHMptWprEedLxU57dRek+j9BTcsXl+WWU/gqCyWjjBlZoVcXo66sV7nSPc71ybo4FMz
5Xct1eZQsD9WnRt1K7C3dN1fVe5dx3lTT5Dxty2VjQlC+Rbo5ZSB3NVIGnqSovW5i+j3rrOe7318
+OgKka5F05XfDzymoBx1w/CwBmmzfJ7UoV0HOaipcHIf2rIja1BaSazgA3APb2RgD54FgYWPEWYr
rk2aXo1Jtk/CNxE+utlhW4UJ1wWqRokwzFSPGSGyaQqOOnkFlBLlQ2/dxBs5PB3KeKCifVt1mzc6
XfsoIO1k2/mo14emPGVmh240PBm19vkuUxsGsI7vP9nNhbD61jkgkRiGSbwWAR3goochH6fDXisX
ksUVnVuqFF8vdnQmgAoK650sskib/ro8j3o1GKSRcHip5Umo+1g6sEj2yNcTr/OyiPxT2K1MiciG
N4dV0YTeW0i/i4A4QWRpor8pLx7c7Y/tnH3ZjTkXpD7praxgzW6B+U5qA4j8m7khqR73eJswXttz
Zt1CrDXut7uUZ4BvKB1sDDNASbMLmzmorKLJ9CVA5HS8fx+alioX+HVZEjiQBb3nv5/AAlMr2y1p
SYStaxBQskK7VxcfUXm98pCkc6psweiO6yx/Ane/NzqBMkG1WLH9XA1oz1g04qbfZakuih89vS1R
FIDcuZX6uQAAqaxJP3xGkKlY9/LVE0zIk5OS6KmUTupSt2TiFPjS1d/qJGGr1h+P7wbTn9PLqm2Q
gNuRwRdVF3vI/4yLtQ9C07FFpo+S8d0vgShRdKe0WNbI4tcEGxUk52c0c9nar+uEonCrg2TVQG6p
AaVYCbBThwr6gVRvRoSybE/C9mHWIsj+V0rvfjdOuLjnnQIX9sLZBP/0ShpS8bf8vt3IcWslHB20
FaTNDE7mX/qSRf/avmuT7cPYt7d5/IHTIzmAYUA+hs2LEH5MfMacV21zodCW39XDEYeW7xrrs9/M
CZ2TEAUvl1YLQylD54y4CYIEf4id/RQCWYRsCbdvb/x82QA5Yf7VsoX39/mMj+E5JGjjofRWgypt
pdcWQbZXVHbIE0qZJ0MgCiT9nPzxNzopKyKtZmrl/UEkVhuXVDN3PgoUoDZpQR/GMvAD+RjpcQ6m
YEHPl+Y1/6vM7Vvdd6VcEcThNy4B1E9160GnHEGN6a3DVPPZkLC3Wb235NzJB9dtJuN0abwwKftR
TKXwZ4EhSwMcnySWUq9pwO3HayHQK+6atG79b0RCU/kczaIk+DvhPLKJvm5ZpoSS5uxl8skHaMWK
ZS1Js/Pit27W1o9gLjKIiTdRAAWhREuJxWyxdWbEroLiztfA9b42WxW4Bd2ja6BytvQuIuK2MX2s
Z1Q+mpYEdarZcIjxoPvPNHmu/lwh1o8kIv/dImyrCkuK1hsYFWFHLC5Fsbs2MJ55i5c+lvKoa5J3
n0q+zYypORQ3LyHjrbB47QXEe6zhFcK0qqx7tAk+ViNnhsU7R3l0iBu9u8PmRlvhaHRmdPMi7Q06
tZC3BhtqrL0PKF507/iTNInTPeC33Pw2PIdWqp+fTAEm9zBKRGTclRKRYq8Oe+EjeOWCDrVMSugO
kHX079QbxDmnKr1aDoPaS+Zj9TElC8eui8zDheYKKH3/vKceOVvlbFk0Cdnf3qAeFlu4x91JT+AC
f7TtObR+3pEurc0j9gZlpkRnta/TLwqTXtaCwW6GnbeX0AWiWyMIHGGdU6TIXgxsnwaRraGvEiWC
7H9f+EXqjYMTnr+fnliuv81fdEf50VPf8KYu+1vIkSZbyuljOlQXdpgoJQj0OzEeNNnDTXh4G3ud
Kk5rQX8ujs/pqxyJCp9jJbPDmwv0S+cYar+f41KKgv9G9AhnXuP1JDas1vak8z2QfT794gIDmeve
vaTVmaWUt7kdzyVkLllUEbi25kqHd1EnBw+vPeeSrNMRKJu8iy0mMhrCxkF8H04g1Fl+R4aP5jfL
U2cEQ0g8YxlflGkBmZo9dl/fTvPXkqPYL62Kgx8+ChRX+HlIWGTheG8XNDYZ8D6lY89kiAjSIyq9
F+lUALTx9rD9tZq65ICfPXDLyzELnuP6VpWM6Mpw5dXsvHg85AJsLC83VCn9vcqdkNhK7O30V4X7
c3KtX2K79LnJ50DxyQ0KZicieUvCQXi2bBYmvxbEqHBsODnlw8kAQof3UhxOF5Of5f6rnw/EX49r
THSFSrSgB86lawidolBRIfqpICEC9YdSdoxq5azDH54gMSrAphdYCVnY4pinglV0ZH6yIToxkoAb
IYFaIncNj1kh8PgqDkOi8kSvVz0MWp8ENgki+qCjgEKKrjrUFEWmodj62PBX1B/fiRP2P9RBCB8p
qZu/V01P2M4JxcFOI88nnZv6powiH9VX4bRUbP2aIm6YOLlHfKwB3KtRnaMA1JjoWxOCq3PlhBeU
X8Ri7skJet5ZuLzDiOb2FXJtxKjl8FSVjv3EBafttrG772c5HBroy6ywo5ZMMg7z/wNU6KpdCELG
DNJqb4xPSsviEFjbqSJ8UENLbY1/kSm7Dzvxd3zn6+cmozIoPcEVIyzvPCV4qEAmJn86eVXARATK
M0Fp4od4x5VTyZCC751OAt5fVuuvWjHJTUkhVW+YChMSEAWaBNgjgg4AZ8YqU7XWdMpVkcpZwl8Q
i/o5Ncr6uiPtB05gNjp7s+3VMDSl8ZpziITzgYJn7LZdeqM3NWDY7fUZOtB8hIaCg+lePmR7IQCk
KmIs62fyBTOkJDPu1TvKv5gW5Nr7p3cIs+wVcfUW/s7gqfa6M/is3eNqAUxNOy8o7sKiQPAXGFxc
IRHzyAkiVCxNepmSvImYN165DxIccFxWiLConrNUFyW1flai90e6pb8DFMJFpeDTkqbUhqPX5tr4
cwr72ukZ/uxCppMEhK6myDpY4wYp8KbZhpiMrLHwzlQGNSDqXiuL8aEWgjZkYxoZyGYP+bYyBecO
3xxYB2ijDmrqcMbWp0tu0XeeEVitbFWizL9+O3zNKOIn/9bR5cJOP2bQ5SyLNkO03ujVt+bMICxu
flgKqCJ2z12T86Ha6J4tDxcwX0ghq15TC753SdVpX0hfWNlcW3ayylj0F++Q3xnWJ29F71DsC8BZ
91ty0D0PVYnb0RTmTGM+TY/vUyNxY+7gK+dFuqPcbKP5tVWVSowrUWA+qI+7uWFGwl3t0XVULm6q
5ROTqINTTjayGrsrWvu5AtwG0V226fPx0magXVaX5O8CRI26FhA90Jp5rkEedWC4BCcI21qySyQ6
mKVM5VFW7XeAmD9FkX21gApEPZugX10rRkPOvQRe9kFN7Cw2d5m4zUWHk+gJcwRPz/kQWkP9sVYY
LP+o5DRydTOtj303LPsaXXrdPmFSjwCOWOH1nAMa2GiXxy7nRfld1fhQqSXzFHimI8VbmvqKrPRx
jAXVTOqiwJ9S34a4+mLc32eDQ/6fi/HXrWqcE+ANAQcn6FHeooSA4vPwDD+B8QDd2kmkTWPlvQv1
Mp5EvcmIv+pcYobCCJXIqx4vkLxHqgr9NPbuWypLSpWC0MCTJPvNGrCDkaoia8S8FSBC9FR6huvU
yHORxL+f1grOO7ramZeszDqTlCO1+et+nL5ncvrgAxcQ1IhmoS9+mhQyapMWvjBhsUrsBnm1sGXJ
NvxbDg61J9K3GE76sZ2DzV4pa87SRmej8KlXpIdKdz3Ec9s8ZU4VtA0AFhr7s9HSlzQM7Nj5jSNd
t7t+qvsD3nEtIQwp1O7w8juWAM7S6d+wZSKQTpXMYlanqJ+WO256vQx70qYGFls7oHfPDf6hALGj
KoJStidbRPHUTK+hqolDg78aWRBBzOX3eFUN6g2wT/28lU9nT7rSbDIarHRppZugsArq1BkF0e8d
64c/GdEJ7q2CivhQAMUk92ReUOtry0PMuAQmfWzsQy9zee0ErrZK6LL3n6mPEEpRhbzLRHusV1s1
8Tiluvic7+q88Yw+PKQxjTjM7C3spYx46fEs354myVWdh+sWZy40sJsN6vszhoJ7HmbWR9eLMXqB
9vOKS/0ZC1QCLmlBs4K4e/CgOaFa7aEWiKSXDu7gpoJd9BTTnewpqQ/71uVmyhuj/eOc5DSj06U7
ukhm26xjoTGnTQa/nnKcZUzCUNtImFpmCk4nosnVlip+wAbYOY62oWFUEW6yxj92Gpjizdn7p7N5
TxgdCGVfbKZqm+3m3/xFOs5WYfQD8VaKqnc2e2fCHt8zsDEYv/kra3OlIHoCXmT2OD2417jnsrXj
Jm9RCTq+O3TA2/dRZZ+nKd0S/xfVN9w55EWZvjAzcnijkkGNnWjCfOwYUSIwF3Ojsx/5DYbVUGAa
Wxq4B90WoddLxGGr8bhM+LAAtOGiE1+g1Atwf4BPO+Iq4szeg7Q5QvaXmJM7/tN3ew5F9dHNmYbB
IGLXCZit00sxyN0DMC++rvCi28dgoNt17z2+KajDCp+EdtpUrVacOWaMJ3R2wgQsxfB0DpcxLKXQ
idoVXKYtktiDETzmt8ePKAkHKnvqzAmc9N+vTmrLfJE6YICBiHWnvC7sij2WVznAltVtzrvMFb9o
hssFU+XFcAew54/QjFooQUwNojPjfGzVT5RbUKJTcUy8PZU2r+aa7ZSIWYp0pFcHK5vbz8F3itwo
BbZUboTRqEa1kT8C3TAfu9JzVNAFSPoXZDHYRF14LCaZV1lrffLrdMngRNtCa5R/zzH7GDfOe2Os
E47yu0YC9LAgOViBJTfPTWpGrb6DYA/clqHRZxx3BV7q9WsnyEk/OTiiXX5hm4o5jEOKLMf5Y1j1
mIELWh1ORkA0gfbz+Xcl9+lsMhAVZeETIdqrykr/mMlK94unVxd4u4rgvy5XXnjM0IP5EUyw3CB7
XBAUz+Zn0q4/X5d8uyFEaU5tNrRWBRaf9pye+qCitQoqkwMubc5HHj8V0qmNmKeeLaz0YWeUbrqF
2i3NOGz6BgR+SA7cB9YJcJY0PD57kAEXPVva8YvdqUBtfLsBmfhlYt/tOhCTZtVUErj7K5r4Lp/N
uKlk2N4/bBsu38sGMvngZdYq6M/yfd2RyTzJBeKzVs/D3vfkkh4IQ1+732rPZAcDBuz9MiKsqRFv
duDfN3dT51Dqxj6RBCuCAlkURyQz2e7RLgKqzi6lBNKRiAKQFKbXj64m9gaIRE8m4Z/abm7pSAKY
Pw+Y+5YBzV5p2tGGYN0i8FyYdXKhpWrcGQ/97fsdohbzfQfIIuHsGoEXxtgl9Q9t0SW/Uvr3q8T2
dDrZvO4tD5XQLBZW/UMawvzEfg2PDRs5fEVZnxEcUv7OTaUxdmgzQRAxgT02Tl2pIDVsL51pVDWd
BO3JvdQRw+66nEpculjgdvwih3/QCqZO9718YhA2eGEbS0TWEh0fvYnGBtpIhHrSUgLSKk2Wjh/d
yEyHkqgHwhTbp9xv+NgoghICtt+vV6Jk5yZl7JI03QnmBdzU5eOMTzZvU8/wyl4ywGn2y/Q6Lf/g
2O6YYNg1TVhYk/9WAEd6o5XvXCQ7nYswdY0fhwIt0MobW3h2CF2U1c0Hrguaf67IShMd8vTEQj+6
g7q9q4x9VqbkkNmwugtGu5p9J0AxIOpGb+isjKt5cVGVkY1bbHH+mJjqVxjzmpPX0PXHSnjWxY7q
dka0ygHFZiVYkuekaFAs1x+vxQM2MxPWkrEYaSqHRrXdQZjlTMl/DuTBvN25wgD8WNbgUsXCq3zD
bv247UZPojC/IPU0Ud6LZDS8hhCaYERlunW2sU9rKeSmrJ1IRu+3SLYxC6zD63azAYyPSBCArpTh
x0lylKnK/FRcHxOmFQHBAcdQ2zhi3OeJWkxFz2/5jmTKTNAq/BWy61vEM+/i5sg/yFuO0qJ+rrya
juD6Wa9o/BZihgRFPRkkKWaftyYDzGddfUHwOkZi3pqpncegkFwMEL63xZd50qOG3GoOoi5agHOP
GqDJm1kD7cFLLqkpyfqGJ4+UDZip2hzgDFE63+QAm5z6sz5h2UzYiIGFVdoLfkt8boXMCrhRqaQK
jLsMk+IELHaGKCkbIDIOMjTRiDMK6daVvQuKAp00POOdou8Nv8U3ihlU9/wZmS/B3+M5cvUG8O4/
6B2nDApUWnDC74jgm1zqcSdSiPh7rvUV1nFtqf4k9w/ORb6tTBnq69TCIFO6XCgROVirDmeYrSjW
5RqucsYUhW9/t/gBRycOVwJgzSbjeiZcQwTzB+s+uw2M3ymwnjiUcW++dNaVfuCGdJCsgvNgO0HB
f8xhTrQ4GiabKPnT3rQIt1ivGtlqkL5rILU67dfGhTMsBlHOD6+hrAkWEUrVZh/GQM/0EXiIDi2s
2FT85c+k3YoLlheO0X1xxqpslpdQu8tic+hDPKtyspJkRJUoEVZadHvE99ywpYYMoD5RKanxTaZZ
eIruAw4pQGGQ+cCdBgoRjxoYRPW8GNx58SnHvblBCVY5paVOC/kC5rTJrzg/mJVNOObGh3yybScp
1bM7xDEfa52a2iVC7I8QfJAb4ZVoDJM04GqsqPyeEcAJFLKMZeSWC69TMl4hEMl00ZkpfCywaEYx
pRbmLXtU7Ei/wsaXnjEvv+Fd4HCDFPDDt9e+0wUMOW/UMnqqLt7ujRLEp1XgXpOAmIOOrEL0erL6
EBL0/WOSXYKQNT9Dwv0mxuhKlK9iK8cWYHwLyAXQdq7TCR3hoS+boR0sxfrTF+e1QlHI1CJ/XqOz
Q4u3R86EvYrm8I46pAWDDpBpvVX64IKl+jIK5pHFPbEDSbt72ZkCUOZF116VJA2FAvgl/ib+Cl85
8mLPA1jMfvdiIlUkanKHulFaVuY+h0X1nAS3sR1dreXjKnnMGRSWHqok61LZPKQsazXSExmY8E38
Z4/FOFGyAk7XAtHLxqfWnYTR+FrqaJN26/I0meqkS2I0kDWljHxj1yaffGDlPkftQ+aCWmJT1D9i
PLYUJbvACrlNsW9kZVPswPSFuCLcvx/Jhl/LpaQxOGtOdu/k5JhkEq6v4b7JiZlxdM3oPOiraCby
La0WxTnEv4olVweNQdjG5j+SfNVrJUNoZQJ7nkXp4UwhcQ2fdAHbl4BDX5d36dL1CY38twHo+03m
2kreCTdk8+3C7U4ME/IFr63c+E5KCt5ojhCQOXSMUF4H+a9cbGLcdkWcNq/3vWb3vKVgZtpdXI83
EvMfB4IKLzoonrzZ1nw6wqb/H8enzkoDayvNjC1yK2IwUNKivub2xFgCTkVf1k7V0qDnyizWD7uQ
ORoCtM04xjiERUMMymgZO5xfSWWT9I+hCuRPWndl2PpliCTBXwNB446hoxwEoByx5mrRXvsasIPf
Zjn53fb3Tqjv2IG9YoAMEt8TV4JtzTYWwi+DNgJhXVo9W2BoEw7wsmJSGajx/DhiR2f0MlGwkgXj
gyVEMFszIGOuJfuBFEA05es2LwLTDjgeEHdFQnVMNp8XJR8C+3Xgl/ptVlYxa4zcPNSVnhe51qMX
oPhgu/yrkRysSKQ6k0H9wlm/bU1GvrAuxT7aqi+zzifAKeuFcjbXW+xQVyVyqgkJl86g7lU9Q596
lznlMzYuyTpxxVvaxUaE8pIoAc2n5UHEiGy5N6Wg+ix+xIwS0QzzfZk07yazmWBtSg/77EVSoWyv
cG2nuIXfO5VDGT4bOemuiUFTKApQU/8XVisON8V3uddozvYaKkGsw4l61r05L3/LB4wbebTvSXx0
0/OGSbsc0A+xiRGK3tBOSwcSI2mr69wWLuCu4wVIsRvd+JCNTolkpVryRekFSSKlPROleZwbm2a5
3Sv/x1pytZnnf3RghzTacntaxytMUtNiL+ofb/ZF4q86vkdKiF7Y9z6RnGV9keOCypSkk8DeYhGx
woF4LKAvzUUVTDiZ4S2pOEOZVU3knBSV2eT5OlJ9emdRBUfGw+YtRn+XUBipaljTWhn22JDGOguW
1+FhjMLNKrpgBbqryp12D8u5LIT1KutVJFWYb/IIknX5ksrvo12Gy6l6wgYos4syZDG0Y9+MJ3KA
RSRtuAlBhDVqNLDxqmZHZdth8GSkIxnWlLaFzBX43AkcozPyyJRuctvL4R+YBnE+lGO21pQP+SRK
v/saBB5/igjj4PUJ9IhzhYaHIddpOWaIq5o5j5mMmFmfRj7JFMOKx/Q2Ju/JHcAt9RWQTiWvxutM
1NF/b3RllekKdyiQvFBb8b3l7N9StePokY2IEYl8f8N1rGVt4MrJug6GoCtcHgHE2Qqa7P0Sagn3
3bWcxfhflb7rJRuLExlUpgyy6xkYY/HGZoLzPiDyWCvCRkq9xDSekjmt2873Tk2iWAzvZ3g+b7ub
MaB6WZhtcMquFrDrSdKwZSDHmdXFRiDZOuhJ+/ddABXXCf+nz3wcRMtvvlP1oNFp3fdNRkS5bBlI
CS/k8panvBHH36id1/IMNA6jaQOqsGLiCacgZ7aFRpUAbVvhiy1mvmy1akgtz3ClA2we+fzSnod5
umCANbyiwKVU1Jrm5CDZJqzFysJ2zxgj+5u+Ibj0uHYEMC9evr1hmzq3xm/i4H+IJhuDFb9mzTvJ
BRwxa9oLrXOzlVcnN8t2bmIBFLMQ7pKBojzwGYFMZMPS3+e7oUUlJbG7Q7FnBKUxITF2iPzN4j1L
Rqb1SHRH/0ILyknkP08NunCusJsF63eIpwdX4CyVplMeVzNSR0yCJhR7PHO0zm++aGikIqw0XVOd
RLomAKfoEQtGgw7gYvLVIAIs12ab7jA+JKArX/ZFtONY4HqeSAst3NfXuXc6mNjQBWAjtyKw95pw
R+hkIhDHtIWFlweMCzwZ/EILJIZxAy/603Kub+fy/XLvr5zlGqP956w4RqpwWc+w8YDuHHQttiaO
QxNTila58bkhUUUPC2RWyoywVyILH6dVXGe5wjBMLTh10X1oRRamjTcYiwDSCWI+xP18FeBWYq53
r/4+hDV6WeIKezlplH5pc3WtxTvHAKNzd+yDd/MklGNOG5AELbkEUY4rtpZQ7nxyPawAMS0+chJf
qkUQK3SgRDcEoIewoju2sdjqnwCNVIyyvm/N0DlhwgCw/0tph+QNYPl16C2+qdtU0Bxp4v78qP3h
2VlDcL2wh4VBTgM/DBTHJsE6flkPK4qLLCCHegL3ZdOff9P8B5ql2sdMiNU4SGAlwGMeY8M+jzbp
jEKI8U17RQ7QL0kUCjAv0mu7JBL8DT6rqE3bk/AyZxlvvjnegAyVxBvxLV3iBk7sh7YBpL+eCcvO
4zJC2ul446ErNhNB3ShrXECR8pNMOn4v05JfMrUn0oDgGZQWpkU2obeNGis/50bPvLprGGd1qGwP
yRBJp2EjzrTHku5s0X1CzKeHgPNkaCsdd/fE6YpyKi5kjVDiWu5LPDrKl57s9rKHwjtGA3knfvow
Quf9BGU8bjy/E6NiuedHr7D2D3gYuSMPfIkVZl5MmYxmTW9jQxbXgk0H0rPzkOUexhL2ZrXAh5AR
L2umLF4iRFvQumiRaDY6x1mrZW+tbW8ZgBkcPvTf3AUW7keXvc8ulRhj0X8rct9AxrYsG4E2PAF3
PXDsT90HbrCHMyrAaxJVQK9QEUpiy3b4u5oX6IdUUD//X+6qqLxQyLKoMOkuvtNbEzWNSTfeydp3
F3Ht1meCVLxUQ6L4PICfwhmi7dKMxSg9JxMM4HobgyVfMas/Ac1dcs+hQlURakElU7EN8xbnFcvK
PrS5cnnlRXqiY/6KvFbJ+cazoKESemQHFMHrqqYCOez77YUZENn71JjnCtxRJ64brbmL0ewADYfQ
bogLr+CuVoWnuvwIHQBcRwaxmB71xyotTsbZMwXtK90il4LIBGCQY8k+fhsbzCa7O4luqWHZZKKG
NO9ajEZzmE5QWEGi61WkqU3x1mOca3zSJfUpgIh9Z0VKMWDrXdjTIFIBL15DLYWb3GpcY68fbJ3z
Tn3sabsESpm9EZ3O0PTIWlSSR9uhh2qkN2hxB+DwOmheJ2g6MpfHiXaY86vYrmiOVCznAFMd8+0b
BAPp9mD8EQlDdmd+2azl35r1X6+RADqPgWZX/wze/sWuybgaRZQCZWMYorRIC3gGlgVMBW8Chbo5
oynyV9j2Gn3BeOBI1O7e0hJFb3G14XuUYUHpEAi99PZShB7YYLkIS82+tKjN17A02kTSUtMrKoGl
FinmcAYfK5m482S9wMcVx9ox86CkHgxLFQoquvytN+j9fzSeiyyR5VGfLL5YacN4l10ueeY1YGlx
FR8WTvbOIYUhxpBdE8CZ1nGhwCvcJc+V31ZsucYOLclX4pw12DEPTbJXndbh/3KyDOTLvigqQ/ri
c0MUo97Eeyyl0P/dShxCcTl00ZwuVxoNROCnnUCCz6HgPfZK9ah5zXxwN/jaHKVe7d2pnrzhVOPy
a+NGXmUogVLLNvzgJWW9WaqPVA8iQIPkYx+v+uxuF0Jf4B5VFdD0bYlRr9WjC0WYAUarho5MKP6T
a+bPvCHR/8GrVrtBdQVGGiFOhbusT1VpybMn0XCPCjBGMzUbgxBzSgCp7fYuzZ2W0bhM1MzxgD9D
AJG/aHpSy0J33OrwCKuVIrYzhc/D1M0pqgHEOv6QfMzoIrK/Gl65rGIVy1aaLi1Lq7Vlcalc6aq1
au+XWy2DT0AvcN2RAqukq7iitluwj0v7pidkHHRqlnhKoBHsl2Xo/v3kh0q3UEkWJF1HMp3eVwnZ
8N6Xq0x5DWvcSkHCZtSm5ueS3wG3gVy87CYlABermpYBrtCjExlH5WsDXLszV15rIek1hss9rTvN
JxVAR+g8miAFLhCaLoWEeNipSc06C7a9cNFy2qDuz1LmGSVxV/ejwfM1VYzc/g8sPGswiW6UZ1/6
t3ATEu9QotJQ7Ueouco4e/luIP2Cf3nx+S/eEkiYLrZ3dRtRH40hQ7/kj6A4lcyEbnvUtQHw7Uzl
r7Zwn48TC8SOOKqgCxljpUuNxxn0iM0IBLlxyF4yiib0jsSdH9ZRYSkpTApR+nDSC1/wLCXB24pX
TJf2mHaGYrAFJYSLIRttG9NGIWASCPc5VGYTTH3QSA79PhWoP1/9a/cVUxYJ/SOwQKzkOXSIFE3j
Y5+dLEV/yvvOxeIKi2X+LBU5Vj41mNjrJMQJOCcm/BeXb1vvkK7KpXOeSWGGCJ+PqBoxd82kkZiK
rDZsnn+cCl2VBXNtJ8y2KSLG47EsUcDtt225a4tIoxE4XoLZ0P9c5SU/XdaKbItMRBX3bQvIfLcP
TP/enjH8a9e6YnCl5aLSx7z9pwis0t5G/75T+Mxqvmhp8z9rMop2fIp201r0lXMENatCZU0/iGG5
O9KKeHIPiasU6W1Mu9KB6kxMefiESpv7yRwORcEQ21jXU7PBVym6DUDTPyHIQgo4Pu6EaxoL1wLn
4LDKMILq7Sv9LauJ6Oz+ee04ftg/Gb7SSVkXrzwVnAI/PzuxzmfJ1z5AZsybIcHXsmTOCDnpzKmv
KevvIJlzvTKS9kbUNrehcguicLSPrIprZktUwDK1wbW/AP1jcijMGwfCllPmeBBrTXgvi/S07tM0
jev4pI3LbL3ATREWA4jj1kXireZTA1+spu799VdDWwje8CmSyOgmiO467HlRv1rKff+3Hqv807PE
nyZvYF4lW1IEdIuE0Dt0MD1krv8G8r+tgJWGV41V+uUvDINLxEQwHspcHfu/ahfkQsi0e72yIv5z
uwyHT9h1xMlmnxyIs0sHhzfci2mWNm7dkL9tgaTfq4v633UZ+3P0k1TTgmOsn+hbxEW3jr8lNMfY
ejtbtz1TpxApKFTTf1pi/0a8PTaNPxyBqOkikc8gsUZNloeEYZDQnK3w3k/57UsTBcZxzgHfjBXl
Ao19+GckvmjGS0WeBdviV9KpK2HvxXBiu3A2kmC+GSANUtY1mmaeoRoyJMyM1Y8WigQNIG56oehs
yMyAhG5sH5FK3BK+5G9rVIMGYpyDfGyzbeOLLaw3hB9p2Dhm88xfO2pDDDdyJ67p8aeeDyrzKBiO
JZiXZdQtZZBx7qshCt42Hy8qeFJY4C3g1ab89GOMRQIgbw5/SUbmTu51DPxaYGmI22Ts3yWjjNux
yL4q6efiPzfgKS0S3EIttLVE+CbVB3M2oEsTaE3j9AR+1LRkvdTd7HLSi9yIhk8N8elQO2eIJcpX
LbTiCIlbuwRKpnmu1bcz6W4Kz3RTDQZ/2ZSNj6zDOzhn7G9da7UYNpjo2zoq7CQgp7+sjsN3gWZs
Z1nhFbXIG1+iDYSmYue/21LSLpWQHxmrEzJN3O2sg9Ha7j4j2/YwxNIZkq/5BE/c1lEyTg1tNPxs
yAfVGfnMzpCmYPw2sR719eH/RqrZJBbo1Y97snC4pumfMMmCklRQeOu/ubs30muikalTRlP2CPcS
pkwymGwvLRAHEdDdoNKf1R9DON8FgZ4JCzl/px9zmRKtQxRSuWNtHeBAx4/8AFWBbd5QoDB/7ZYB
dL4j+rG2vSMJxHgKcGwZYuDw03Ww8FxUL312iVbPVBf5t5yCnDwv2YkxjVingNpze9ZvhTmnuTBl
/w7YL1bDpdWo3VKDJ6KRaXuMB4shK8zB/d5iYgeLenWXCkAF7qmBfS5mJhdtyvdRPSSQIYK6+BFl
Wbf/oiXgCsqajd/DRZ1i+Y4mtpTowBwnKoqqFmYX9mQgkCati0NBhjqNmQkBEeOD4rQ0wQcMNAt2
8NepVcwlvkRjDsMZVcTIygzD/6ZAG5y0NE6ooc6/i4460y5SZ61mDJc=
`protect end_protected
