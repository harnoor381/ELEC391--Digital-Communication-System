��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����,�1	�)��&��(��H����dP7ɨ���:��0����,�6m���Ib� ��JK�yUh^��9���E`���K�
��Q/��V��T�"���-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_d
�t!���N�S��گ/�TNM{�C�5���M��;����L�S�:�{���\p<��)�0W��B�R<Qt��Ԁj,3Ӂ�v��`s�HW��眣�U�Z.͓k���ŏ�^�sGt��P3U����ŷ��T�'~�*9Hډ���:Y�����%MJ�I���a8�0�=���6��nOsy�����b�	B��Lj#3Bq���Վ���ۀ$�>NG�K�'g,lץ�E5��SI���'/�/���7��o��5g�2��g6IUN;q������Ӆ3R9�W?�F�LR�但�
#r��+Br�Gj�M�H%d��1[ �w��'��&o�-kh
��w�|Jo��������sJ3s��N]\�+-)k���DS73����#�1��I���_p.��a�Ð,�՞�˗�v�n�[��Rۍl#�Z=�TSc��ޥH��^s2�XbQ I(��/�P=[�ծ��][7�	����9QdZHH����^�"3Q�˜��f��z��"�HQ�n+2���f\1$f��*�I;e��0	����M��T�>K�d�Ñ �,���0o`�U��n���
����Ch�ql5u�'+�O�qխ��:O���WW���@R�S���'�Y�[�^��R{�D�����P���UE�؊�L� ���@٨���d��B�O�h��$�.��]�Z��VI��</ŏ�ٯ��	O�&���rϤ�Pƿ|�Z�l��H�YBp�� "�����luZ�UI�8zv2��u"c���0D���cd�<����N��)�a�p����^�Z����Q�B�����Q�}�k�>�9�ԸT��PA��6�P&��w�+��E!�Yq�Uh���9<��Wj�bvϫ�O4v��MJYzx��������6�:)�B�"ʩL�]�U�����H��V�u�����x��.�;Y����ݳ��o>��"�Uc�Z*�c���b�ˢ&w���b�&��$\���-+	|�3�Zh8�0UܣC'I��@��^�P?	*5�1������H��.f�&[�$�(��޿~����0|�0�s +Z�~��G@�P��#V�Yͥ�gmNsL�1�!��_;	K|��un�}y��Z+!�9;l����#�z��b6����肘Uo�%
�l�k��ٳZϷ8#\� �aV�z�>�|�#�1��o�(�x�0�/��ub�ɟ@�µ���\��v"2���'���Aq]���U�0�?�q�ـl��ͨAy{DP�zmF��>��L�fy��q��\9IQ2�W�M+��|���Ed'���2�"�L��L�0�J�<-�ח����nC�8F�
��"��A�9JgH*y	y��*q1��]G��S�4�1����y��{���
�m�iTxl�Ir���9����*�^s���H��e�骊Ү�	�c���m��|��1�G�KA(������˫iB}��b�[�zܴ?wP� @��	A�vg��3y��w�j�Sї�}FM~sl�b�}�r.I
���y�vq�p��|��H�	��m/���*n1���!_.�� jj^�iEï�к83���A5��g�p���C3���������R�u}5of擓����3�X]ܡ����B�S%nī���6Cr[�-�星��5�K�M�2�ˎ������~/�}�����0�C��yi�u
!y�r2x�Y��ʜ�����3`UT�m+���Nƹ����C�]<���O�4����ˈD+K[α�H�`G�~A�^�j��j�G�a�6*��TW��Fĳ.�2�+�7G�Aq��|!�mv��F��v�\'�/�S[lL�p��7eR8.�P/�S���
\�e?�/�Y�`�+ۜ��BUC\�l[m�6��??�G��++�"����e)w��5MuH�:p�_���WI-$C8�	 i6N��q�)a^ۈ͝Lנ��-�5Qщcs�\��,)y+�x��H�ߡ���X;U�ξ���^Ype;˰u����ƹ������
E���a~�[=�?�*�^"]D��߸�B)�s�Y�l';8T��g��P�3�H��ʟ�R�o��D����U-�J��UP:sw/RO����YS��p !�����B�-J����L,A@���MS�r�A�r��MS?g�7���������n[�&�-jл��bMV����Tn�VJ� ���-6<myU��~��?t���)@K6�!�bY���b"��CT��P�N�H��u��U�N��PK� �x0K�'���㘑��s��i$�x�^��im�e,�K� J�H�eJ�V�o!ٯ%��N5���	F�����$��ͅ��-MPrh��%-�o�v�z��%��)3�̬*�0�?F�4��a>Ǻ�q��ܺ˞M������c��v��q4�Z������@��g&[���a��|�6j�]�8@��/�G��Ay}��_�����ʒ>�ܒ�I�C	A�`�E{�O��r�	Mt�zn/+�;)�#�(��ޭ)Β��W�j���㺠e������������j�O�6}��ЪM�U/M��~נ��ꌄ����e��KW�!U<��bd�?����O䓓�" N�5[f�e$D'��?�TB�#!d��\ g���ٹ���`ZZ̺_,�1=�i˰F�ɸG�loĔk7�n�{*r�F,���J�l������%zŌ��kT�>�� ���N$�Wi�9;�.�4j$М^^��E�*RwoB�B�r�s�TZ�����"��������o�2���tj�ټ8n-�]�DI������!I�Jŉ���A�_l��39e7'�Ch�ڶ�ȴ��(5���>X�,X1���|r����o�&c��B��� �-�� ��:�8�IӮRkc��6�fI|��@擪kk1�>�2�N���:��ј#x�o�]mĩR9o ��I ������%�R�`�sE7�T�ͅ�y�b�,v:VS�N\ ;�AVڮ�~6{��eJ5�SM8D��uFrq���<l��Yw�=����e6�ԝe���~O��[�½!]�FU�����@��{��$��	�<��v��'������T.l���+(
�}�OĽ�֐-a�!��G)x:��%I=,���9�W�'�R��͏t�~�!��Ӳ��?��&�_��S
�՝���1	�HІ��H@�d����_k�S��6�ɽ$a�J5sP�|���#�6�&\�UH��#��V���(m͢��vQ������_�-���w\�z����?��O7�.7��b�tb���և*�[�,��
��Nx&�x�pH�)<k�뉜���,�(R��V�>�&(��~s!����k%���/!1��F���*�+����%Q���_�L%'�[���������3���[�CN��/��8�%���ɞ`����\�"
dL�fPH D�:����j�l���|��-��*�ҋ�M��A5�8�\I}
���h�L����뼙v�F�z��>�����s;bϬ�L��mӅSuH"��f����+�����fwO�v�m��Λ���� V_ӊ���YE����%��Bc�;��8ޢ�\�3R����b2$D�������� �s�Q@�8fO�c��*�m�ּ�n�:�%�|�q�)?�� ��D]��@�8�<x���xCa��u�2��C��i�y��P%��i� ܩI��-g9��`Rb���= 7�Sb�F�{xY�7h�p-2v�֪Ѯ ��λ�Hس�6�2L�~"W�$Ψ���Q��F���Z���HC���1��<���sX�#�ts~Iy�DgMut|��Z�;Y3�,%<|�*n��Io�<��g-LM�d��a���e�*�gw,_�X��qMD�����7eG���|�'=�@�wDU4ej�Ь���>y�C�Z�z85(!3��S$��C�D�7��vQ}�p��Wj���7����Hn��Vv��"�Oa��QZ+�[PS�'�u�(�m�H�d���;<�8�u��?�O�ш�ĉ�}�C���'Av�XE7^��:?Un����Iv�'�w���]� ��p�LP��,ߨ�@���E����@��(P���g���>��M�Uo�+���U�&�vL�Q$?����Nu�F�XJM����uu�;rՎ.�8~ �g���������28��E�
>�4f�R�%y��ۑ��9B���Xk�ٞ(#�5�H���Ɵ)g���,��+�����/��G<�J�;��g���X�(����{�,T�wl��,k�!G�����A�t�b/�%�J'<X@�t���L�L��8��wA�.h�)����3��*�<�71�okh�kewUm���_�]w�C�/���7���4���S/�A����P]�=}��q����rjy3U�u��5��wSL.�����z��~K{o^��֌p"�&��_y�".YV�M���ƳиgD}�E%&J�N#��N���I,$�Q�*�^ <���<��!X��vl�J͏js�z�G�b�K~�Ɵ�	Ȑ8��M�|��Th$����u����:W��`���}�_ł��<B����Xe?Bd
5���\�2�=����p�6�Ɖ
1�O���=wl8���Ej��mQ���@vX��0a����X	/D��//��Z	�)<�[�\k�h��%Q�<�bƬ�X#B������i6j^oyL"Bqԓ��%_��k�"��S6�͋f萊�̒�)}Ew�Dz��՝����\7�N&��Q�}^P��[)1�����#Kژ�E���A���֚����@Eө���s�#yE�&=��g?���/t��c�;����G]M~���l���f�*�����BX�� F{Ъu�{��`�H©�N��'���:�:U8C'��ٸ������ȍ�Ib*�_�F��{�ʺ�p���mS��N�a;*1 Ee�K�Du=E�C���Q}!u[�f�8�J:� <36� ��(��F��x� �b�̰��H�f���C~�C��>����V/�z>�����h�n��QFc M�a<Y`�E��2��y*��/Q����xR�+hϞ�uަ��Lp�v�y��4�)'�8#�h��w���A���q͏�0����ך�ܷ���b���������wx�#5�O�T�a)D�Scҽ+'�(&�j���	=�!1��Cx��
��>~P�p�p�p΄��B/O�ܾfzBM�t�@+��zrn��W���6�)G�M�[��~p��%i��H�d�͙(ˡm8n��n8�e�Żoj���f��� p���gJ�Lz�'���Y�O���A�v����F$��T�?P'�4z��%_�u�Ƽ��p�	]��>�d�a�r�Jz��R����#<`�
��1��$�O\��O8�7B���["�\�	u�:UJغ6	w�$v����A�bm��� �55̦?Lֹ��K���H�O��}�P�B+3�xr�0Z8J����h�ƒ'S]���������V����0��㎧8�1+�忼�N�*�C�� ��(@[�����Fsi�b���7/ZB�s��S���>�l6�����i�X�q}�oX��?_t[�:bb��+���:�	��>�V�}>�B�����5`[h�_�梾 ��ї�U�nLs��W���m�7ak꠻�.$E[�y��a�r�T5~_����qc *׆������8�X�:2r�9P||���"��<젡�Au�_�����2�)۬�Z=뮍s�?C��T�%2�8��n�y ���؈�P�����U�w���'����4�v ?]BK��E׿��e�s�)ϣ�B 9�B��_�1�Mw�x�z�EȊ��,EK1����{Mx?�
E�e��\q�9��u_��z/�3���6�g��λ����IrL;91d���8R)�R�q?)u]u�2f����#q�����.3q0�8�h� ��ԙ�;�������1x�S�Ye�<8P�X�L/������?���	B>��:j)ּ�j���q�����:{ʸ鹲>.����Hp���x���R2��oS�-1�P�������SP-��r�?�|�i��]���D����%�t9��I7�vMp?L/!yP�/�͕���{#��Eu$�\#�5��Ev�6������!�F�)��aϴ��]�|@�{G	c1�־*��^�<6������[��俱�aU�N�E��o�ј0��V� ��3���C/a鯮<�����66��A�'�Q�P��9�s��a�:̅HE�ټ���<�;bU�G�hf=�	��+��� ��b��1�>����!�f;=E3����"A��,��s�nd���[t��9j+%�����P�[ A������o[���+*HW� �?¿Sp�>���g/�5<�^b�\�11vt�t=6*�&.P�y�l\����TJ��J��.�y-��/�zt��/`d��L���'���Tу��Z�����m:���b�lKň3F�#H��$'�<�d��U���X,�:��ӟ��ww���9J>6���^����Ai7������Թ#�t'���1��c��M��[��[j��Elޕ -y�t@����>x�\�N��L*�^Ofٞ+}	�J�y��q0�y�ʧM5F}�i��*�D�@h_�������SLx䨊'�/���	���r�S�4Z>L�zrѠ����e7�Ax'Ch�P_x�����P�!����F�ɾTd���j��w_�=�-�]DDN���|8#y9�x���I����P$,� �S\��/CY{cAgP}@�HC[ �]��]©�l'Y��Y8���4�	��k��u���w`��=Ͳ�
rڷ�nA��D��C&m)i�90g3Q��?(�G�;8��'��=��vq�����Nu�hKGX:���t�����$ � `�Lȋ�h�`&0�ݴ)��D]�W�^��ߺ��h|��m�?��װ��l�5`L���O�5��A�R�⇟�0�o޶��c.wj��҃���v�s�C��ȽQ/���{�"�v��ȏ �JV��
�ҼuJ��L�cfm�۟*6��V¥V�Ƞ��i�s	]��q� ����J<"P��5��Ƹ�q�a5�}��a��F���[�L��2YU63�y"o�@AO��C�\>˫/��� AS���I�ֽ���°I+S���LY+��A�oX��/�ʨ�l�|I3�+�����:^���]������X���S�h�c@_
k$�ש�+=+�f�"�?�H����5�~��U�G	��$g Y��{��GO�c�FC����;� %�����2�!U����/�.��_4��Z�`yW� Ͼz(����H-4�)�g�`��$��׵J�'*A�g��/�Fa���
bC��aGvy^���8B���g�u&_v)!>�ʥB�u(�ID��\W���kOy@�
T�b%jT8�;N� ���|�I��,k��xO���J�)5A܉����B ��Ą?�eQ�t�GO1bG��0�N(d����}8�M�ڛVM)���C��c����8�t�a�O-eY��<���W̭�G�Qg�� ش@y�̐U%}^�\��	3l1<bƁЄ�E�.��B����eȡ���K��S������+?C>`�O��6��miO���ǐ�hn��	�A3�(��9Z��~ja���'7�,�zmgޯ�n��P�������f�{z�u�����5n�k�=\)��"p�Eە1l7��u� 0 n�&��cȃ��47�?�s;}�.��e�����R˷ȓS��Eݓ�|��]*���c���ː�d75%
���b��u&/(���0�)���+��ҁ桁���4�����G�b�;���l]Δ��u1Ј�&\�����Ҹ���Q�ѭ���KMh'$(O�����3���(��C2Lp�	���8����~�F��k�z��e�O��=�!���l�����+<ٕ񨦙��z�h���pc�EU^��2p�=?�/HFt���HE�
�l�y�@������y�̥C7�}謢]S�l[o��>ь��u7I�j�M0�E�\�8'�O��s'j�����5�-[���U&T�_�5^9 ��\�W�� .���))n>>�"�Lewdc�-���P����<r��T�\	�zH|"u[�E^�=��~ؐy<ln��Lw������Ö�}�'���I���}�d����BH��aU����_�l��B�'xO� P�o@eY-mӃ�;KZ��ecu�`t�D����|B��W��������+�������\5� ���y�o#�R����|IzNi%�iiA���l�5i��q/�ַ�	&#9`4�k��}�0Q����T��D�Kj�����`��1�i�5O!2D�]�0_�a]�BJ`-qzk&;,���^���LP��y����r}>G�sq����?��������L��3�.�sL��W��@I���Hɯ����x��P�Ã�S���H��H��V�K��P�.�
#�!7s� ��kw�S��*���2��rc���_g���a��	V�sfZ�a��*c�}%�6�t���1�t��|��)�R���}����uS"kz`���|��"���l�M���e�].W�*���w��N���b�{�W���T��8y%��N�w��k�ѧc?鍲���>�,�_�ԛT�_qM	�a�C��K�q���}Ceju���UE��F���,ǖ�*:6i2'�
+^��safꧬ���)�.��W��P�����'T<��C�ܘ)�釚�[�{�s�4�?"��fй�wz�ר����w�� �NƀB˾��!�S��������K�;�7鯬�Ì[H�i��x�n�L;�PIp�U.x�|Л��H�У�ߡX�K}*�@���q�Z���6f�[ p�d_v���F�=�ȥ�T��z9q3c�1`�a��A)X�SL���$H�����AqͅW�q	� ����p��lt.��c�6T�8"��8�yPo v;�GZ�܊1V9��o�$�6��#��5)H�s5(�W-p<�/��#��Kf�6����`}A��h�Wx3��%�.$����Y�w-h��`�Q:���d��%���Cx]��6�1���C���� �9����W.�|VI.Jڌ�`�~���M�������X�L���K�Z�F�xv/�t,)�'�3���܋q��:�<�qp�Y�"�-!�V��t�n��O��[�xY�I�w����)
���`�H?�-�*��%��$E(�χ#R �2�\�e�M�r�ᮎ�B�YR\�G�3ղeU�u��{�0�K�v����@e{A�s����H	A��|��r#5�4l�up�z���:�?���+�!�C��}�BdA�84bpY/�b�*JIy��#�Pec+bG�j
>�����n�80-�d�s�[��a�s��1��B�|�%6`�x�o��dX���5).�]jx�9��V:��o�>Z�F�P
�M�R��M���24rp�BK,�ӟ��M��6	���*<�s����rT^�{�~s�Ĕ͟�$J�V�m�Wq1�#�XD�%���s�Iԇn��ڣgWD�+ȸzhҩ��T�aLDO$\h�#x�/1p 6<���C)�Z��(�Lj����FIG����RwokX�ަG�,�;���ai���7x�v��y�����S�k]�l�E�4��X�jP�$��$���xY�Uur��H��3�L�p>t��<�3�j�x�����a/ѳ�y��� [�tX��-�c�3 ���tr� ß�*~�@�fI������'�N�m���ԖvV�~,���Uӈ2����4	������mJŢm�8�"�է>с�H�~=��)�7��kc��x,W����c�J��OK�j�^��Q�@fX8p�c���&In���3�r�*�	�V?��Go�����nj[:f&��?������+�J���g��K)R�IfԱ�q2�~�k�X�E"l�v�hctNUԂ66R�l���� ��_�m%IB�b�pهQQ�W��b�Ώs~�4~.6��4I�X��J�U�(ƀ�l�sr�o��Q�U��_G���s�mB�%�z�]�Z�ܞ���=���h9��8�a�xX�F�g����-:u6� ��Xb�g�M*Ư�y��¶�BG,���ɚlE�����޵��c�w�X������=�RF�����]I3)�>�gt-�#L���n�|l���<"/X��M���6���fF*M� �TD�_W���֣�B��Ό�R�;��h�g�r)���HwD-1�3�&���2�1�\S�z��Y�Osr�=�8il��^)������͞X��L���)	B{�fRHM�m�!��lM�J�N������K��1^X\μ
 { ,G;Ʌ���鍛x^���]5�	��H�3�>;��B�Տ)�વW���֞��2Af+��y|�lb�_�,r��^j!���_�n�K��u���I�F����>�N����f��*���|q���_��YI-E�z��#ޕ��"#�,K%}����S��.Հ������̤�W���?9��A��y\!����N�ԑ�j���'�6:  ���xt(~�-��Ӡ�߂ܕ$�1L���Rv��I�����c�+оI9NK*ç�e��7Tڢ��L4(P����ܸ�2���n��d^�'�ٵ5���H\��=ez_����0Fr�����n5EvL]0`�F�q���q�*��8%nT(�Q�0��{�u%���Q
ɥ�:�ݑ"��Yb�%���9's>�A��Q��p��1g:/���S�_2(�e��)���&]���ǆv�VM
TC�8�㤌�B>�$�l�p|t���y_��}C�[�������m׳��:_g:g�ձ���͟�QSc���>o�S����U[$��B����T��ި6�Ќ��C|�B�ރH�3���-�M�@�C�ܓ_;�QM'i��ب1�~���]_	܅PoTn��`3��G{��
�#c]�b��d�6B�B�BO�f;P�^u�іo�C%i����� ��~�q��\2�py���hR���b mվHf���V ��éZ(�;�a�Ι�T�MVS:������O�	�n�˳�3@6�W	d���7��nl4>��~�XA�)y�Z�k��/����}��xn�S��e�b�� :�z?W��㏁��T��k�[��Y6x����~�@��A$(|��L��,��_}A�j�����t����}�s1����L��(S幌F��.���� 3jBd�	��{ q@�����+ͱ��mJM>cp�F���+�����ޛ"Vp&5h}��/�z��ϓ��������ʰ�"�l��������F�4e�h���>\����'`�sv�M����c?VvLa3�e�=G��B10��F�d���J�xP�	�HU���ML"{ԹS��ĬE��"Sؼ�3��b���V�C��6]Uj�g�������=�o����#��7{����h	eb�k�����l�m,��TMt1,�a�q_	�,Y��96�gw*�""��ˍJ)\�D�r��I&�Sg�ߺ�`���]��5µt�k|׮1X4�PU�В�xN~z�v:G9~���x[�L��T0�� &��q�V�Y��!���o��������9��1v�?�D����7$b7H��ç�S�l�)�c�e�z�eA��?���/�@��ld0ӢV=����q:�r�d�+�7���Yǎ��:Y-;L��� iS	��|DL�$1n.���!:4�z�p
i�'�k�xk)�꬈�xz�-Rޣ�����F�^t@&~cFr�'��*M��c��"�$E~�A�=(���ر����8=cy- �����3E�@��L���͢��|6�Yu~VR�g��>�TLN��9U����Aj3��J[�Ĩ�7n�&q�����fO>�q��@K��a��.����CU�zeҦ��g#��G�у�r�V�AΟW����`ї�	7��L�<rߡ��b�����
�B�!Mp�g0�Ƀ�D��ٸ��+CiXX�d4HR��:|�h���BoFұLC�9�&�m��/m߿+rY�W/휨a�����)�2���ʫ#.:lTWpP�3��D����v�H�ྛp� ��h��E}�_�W��Ԓ��rs���J>$�#�^sw�B���������{3Q����s+�6ٸ*�7)�0����ۖ����kCM�R��`�Ei��Q���e�
(�D�����f(�/��[Y뇘��F8�p����\/9$Pc-t�w�ࠒ�=��)�*���mH�#����Ʊy�?2�Mx�YIk	ƈ�lE��PXA;5u�Ǆ*=�Z'w�O7�K=�Za��6�&��~h������]�qI�`�B������)��'���� ��m.?>��Ę�����?���w�I��k�����ee�V?� ��
`�@d�*\% �)-(&�H,�3�-4k_5�_�;+`��F0����Qt��~dQ�S�AD�B
1��}[t��n�v	����|ed��6����=���{؎D00��oYY'Tcw��'�b;���R���}:��*��k���W�}�g�t̩��j���}Z8��0�44T^�-w��s��#�-ga@3��j�1��s[���<���ѩiP~��u�l���� ��}����Cv��DkZ�;J�H�k�^�7�o:|��c�$$�_Tz %�;��"�Qb�l���}I��+)����V�IZ�sՀ_��@�8Mg�Q���Gۻ�P�n֠�F�o|�	�aB�r{>a��7�����173er�t�P�7i[���)r�J�
��Z~eK�M(�^��Ɇ��jN3�Ã�3hh)U�2�ʘ5A3�8Ͱ��B}\�6��"#_�p����Wo����ͤ����QR��?��M��	�T9+i�5��Y~�v����P�:,��Z۶Vy�V��k;d��(�Y%��Q�p������EV�6>���g�	s�`��t�w��i4,�e;�h�)�^����:N��w}�/��e��#;������F8L�7Sx�V���`����\�s\9�4��rQIdꊖ���
+��G�2���Y�~v�of��Z�~M��iՍ6��}M<,٥��b$�]�~�>�6I�'�Yz9�"����_Qq˽=�=&��Y�tw�f��3�����X�7� Ũ<�]$�5��{PiɊ/-v`��]��*",'���Bk��F1-��g�sD{�B>��߮4��b8\K}+J�☋`#(0�[Re����g� �a[(�-l��R�'�|1�e������3��ץ۸�LM�$VS4�!�XӰ�z��GS5���X�x�]��f��y������Eҝb?Jq6	�0]X���9��̘���x�e�!��y��k�ԛ����2��'E�}T0Pt#q\yb���w�"�Zш�]:����%��*i�*Tۉ����<���lM�4� ?^��O��`���0��'�ZI8ȼ27�?D+Y���w�!`��c��ca�SF��y�� |��7+o�QZ���ښ{���Nn�|���_l�+B��@������y>x�u�S�i��ѩ�)�g/�	��0�{��,NL�毜e�oԧ`*䴔s�8W�Ω�t�9��f�M�Ф�b���|�#~®Afp'k��Y-H{��-1.�8�m���(g�b�!��㥜����f�l6&LG�}#�Z�g8_�����Јfj�<T6?ం.�ݨm�w,��Gt���Uq��c2�e^6�^Zz��@�:ĿVky���y	��G�ea���Iׄf���}{g���,�=WO�&)b�(�(�(`0�G��b 9a2�k5�?�����%��]��*��>���<����>L +�TI�7��#��e Q��4V��|'ӕ�qt�Yg�	��P��>
������"$��Q��V_��@x��.���ՙ&�������G��MG�+��6H}��j�rE�r;@1�~P������h�w�qo�n�*�f*z;c@2�lܣZ����'��:���DBJ��=a���?��y���m�����C�n�%$��s��� �A;�Q�f�}eq����ۇζi��3�]�������@��S(�˃�.�����'6?Z��-}��`)��,u/���� PD��It�u��^c����Sݹ˩��7�*�t����=s��~�}`�ژ���ƕ����w�H�"��h,��L�C_0����x6 ���gp���������C��6�Sp�	�qf�z'�����Ҫ�n�*S���)|���v�E���uX�w gi��DC��|dXtjO�<��25`�OcYU^[	��u�7&���K:��]4
��4�#?|נe��0�(�Q�*Fv)��UMx�ފ�H�X��-�E;;F�`e3k���p�(�L���4�xe��9�8�]�y���@�;�]���Y�2�I}v�Rn�`b��8��nU��?s| �H���p�}�
`+E�Ͻ]���VP�8�0���:�x�������(�$cg�u�$�,�7���:�����H�C;2׶��E	3�-�-��i�n,���ps֠�[a�U��QB{W����>�p�B�˄���7��b�͝���^<,�.Fj��4�;�,`��c� ��X��{d>h��Y#l�Ʒ`���%��ѓ�N��VS�u�H���I�w���n�:�8v7�x�0��7|��fr$�h�Wݹ�~2>��AU�1�ʔ�o�m�`P��MPY���U�`o��y�BB�G��L��(��Qy0��M���&r��r�{��Z�IK�Yծ�t�yYo�R�5��su�<#���A����_+7l E���BH�U�9&�<䪒���Rū�\%���ӷ����7j|��K�c3��&Uĳ��8s���Uo)��p��>��*�&wbj����m���!�!�M�I�}�q'4'8[\N��6	t��_��G�D��Q�Ar�u�'�s>k�x+[��7O���6������k�NV��<��}]�p�s ��|�xנ��|4�\�Q�ҟ�D��a��ײ�Ku�-��͐E.�A��DS��b�B܌��>�,X$� �mf�#^�g��'�ĩ�l���_�M��l��>��¦�V&�`����\$�8���~�]M��������̀�����P�0k�rH��I�6��;X%UH�3����3�v�����[��v���_V\�O9����#,������A������(�4ù��}D�H���q�c�|gij���:C�I6^�\�n�7s�`������::��(��R>��f�������-~��ME�A �X�'� j5�mS~����@!��%cm�G�
�[i���,����;�͜i�V��@Ǵ8w�~M��`�~�1�u?�bd����~Y5�t���A	9�D�����t�C�R�����F.�l�� ggV��X�#D�C���y��� ���'(ݵ�N4L76��~�|�C͸��죉���VK0r�KQY*�R2��kt&W� <�\��E2?�� ����ׅ$X�tVq�ö\�����3�~��˗Y�t�iz�ul�]��jf�?�%y���'!������3� �;��o��AȞ�w� �-:3�p�;�����&����)T��ey�#�&�!��,QS��:��qat?���?_86��@y�<�.����T/'󷤓!��i������DU!5�RW{ؕϸ3r�v�����_6��ɸ�J�Z��FdЀcқ�i�1s�&#1Cٓ�#����q��3.m�d� 
��}����V�:d���Ϊ+9>��ҥg�I@�N�E���#})���/W�j	��c�j��`�j�)�ٚ0|������@�עLv�E�ȥ|B����#n<��P�o�C-#��(��Z�d���A��7E����t�9�+��K�������V(a��S�a��'�R2RI�,���5�c/$H�� ��p���n�<�6�dY6��3��V���]D��il6�7������N��`�� y9�0�+����>����~v���Z����Њ't�������qݟ���$��� @���4�~/~��W���LvG*/�APE���J<�	g��������C���4c7��̕q|�����se�j l�7r^X�^���W��AХ��k:0&#�c� 59�H�s���@�z�"�����JKբ1޳��l�'�>
:Eb_��;7�wg���*�B!)�^����M�Y{�G��~�»��#��`��O1C�
���#~(���Ё�Ƽ�,���B��� �b#n]���*Q����&�p�+��J��^+k_��w�-����2��gEF�ν��|~�I�����g��+�L��:?�M\a�P-�ɩD�ˉe>,�}q�.��1����Z�AA\��!���tqݼ�D$4��Ph�%��'�����j	�ԉJeu� I 1���s��s�t���f7B�߂���U�I$:w��?HnP�|���l��g��_�#���qF��@���wZ��K: ���z�z`%>c�#��x��A,�!9���M5E�鳈Z��-CA|¢�ĕ21T7�p=���p��h_�	E0��� ��v���CS2-����)yA��&�=똶�חF�o��Ƙf���X���9£,Mli��� =߹��l:S�".�ΌkD��ܔ�4���n	��@nW�K�xP ���ت�P@�:�ɩ�+�e�]w*��|E;����3V=s�b^�������ń3��!h����i��Ô�ςJ����Mg0$ć�
���!�Ejq��$� ]m��_L��o��?��Q-
tn��>U��}z�G����zE��aH��������C��7f,��$�����s�^P!�e/텐񺂐S��@��_F",�Δ�8��(�� ��� V;�`x1��$&�>�%����Rp
����v�v�I=_IȞ)Lh�G�ަ��vd�u�<FS0��PN��S���R�n5o�o�2:���%F'���ߵ�v�˂��?��|�%�?��-��9R��QP2=�k��d��2�CNL �CZ�	?��~M?�&�l*�tՀ�� �@�Rxb\F=���N��'3Ė�t�q��*BKs*�9Z��9fA.�* 4n�����P���ʖ�5*u��`^���:z�a)�ɽ#��B�:�V�K,�=��f��j�Y�^V�Tx�fwu ^�kN�A��2zt/[���u)�
7e1�L��uN�n�BA���g�<}�uVd���;�����X�`��
�5�-u�F��_]0��vϛa%:s��{�u�gd�3���&���b�t�F�=o��:;�<P�Ԁ,.����i�<"��:���^�#X������=71%ݓ�Ne~!�^��2q�%�i P���ް���b!�_�ֈ��!!f{k�x5����%Z���Rֆ�6f<�3&r�Q+���d�D`��k0:X=����a�>Ɨ��c��
ztC�GZ��%�O̯���7;��*&����� ���c~�-Y�X�e���f ����C�\��[-�����w��R��u�j��n��Z'꿴8~C� FP����3�{AO�+��8�iX����e8A�!r~��y��l.�SN��1388#��ۺժ��Tz x�On����Rȯimg�+��c�i2L�J���\Ԫӿ�WC�����;~s0<~�>q����e�n!!h���G������	b tD�7�Բ�e=H���I+�����N���k��[0�)@WOSP�2�Xq��e����:�V�	�ȩ��|���,6����B�ٓ��E�N� �B7ըmT'{�2gD4�Z�̿�=�K��gq����I��n�e:!�U#d	#��Dt�R���m�${M^�B�Y8�J��T�81�G�fM}���.�
��^c�m�e��/T/�� 2��3��Uo��^��)av"-Y[(�oDI?S�B>��B�#��xzk� +��B4	-T�>���m\���D������Ulۥ�٫l�|@���پ�Y_����^zx����#��|����*�_RW@��Yf=$�������Y���i$Ϊ�s�2��9}����V6�壸� ��� ;�L)v���ޝ�O%��Wq=#("	�xd̓b
 �c��ks&SJͥ��ڴ� �j�jx��|R�C�c���*��'ү׾�`鄒�/E]3�x�+:��H�"�j��GC,����8�A�|*k9+�Ts���l�"[[�&��FuO�cpR�s�m��	nLym��1���Q f�Ь\��������	�OL�߻&���������Rw�7�pWF7>��{�� �LQ������"�Ƭ��r���rA����4�Y]�S2�n2����wA��_Y�)D$1��&J��Yw�T/��8	��4*�r2JN@�:��P�5�[cѺ�B�+޵�}�e�����o�~�P(�|�>����S�1��p3+	o6?�sB�s�q��9���A8�����KY�k���@�m��i����V�QE6v��I��'F�ZTYg�[��o$B)����.O.P����#l���Z_!���͛�:����am�B����Q����Ѽ=�5�p[�WY�q�rK�Z"�?;���	�vs�}��?�&���3v�sӂ��R��>�MS9��/
}jق���,+�B�I(�v�U�/	b�O�c�T,-��1�s%��HS�X�������8Y�mZ�+R��)9N�˸���N�m[2r�6�F�����$i�o�4�<R�X�j��m0��t�#�i���\���@��r3�$�Bu��X�
��ɎҘ�g���Y̴ZGVYۺ� !��*�ɲxn�3��z@�|�L&��@;C��`Ř��q�Z��x]ˌQP	��i���"�gfd������1����ܕwm��j������<��`I$���༰S-��7�r�!j6䮅�c���&�g82�D[G�����C��7��n�����Q �ع���WwC(�q�b-#��2X$�o��U���s�?����O�h�Q��-*�[����mB-:��͟ԅ�E{M~B��k��J�	�юq��mĲ��z{r�;�v��ŕ�~�t�4�V��hf?|��0����{s��/�P�G�Q�-�w,{�Qڸ�����<h��T��i+deWR�Ke���T��1�M6��J?R2���n:����P�{q�ޫ������f�9�<��r���(� [W\��`��&�^0�[0NތB`�A;8U	�0~���;�4�.�����fk��v%H�
wa��}f�pNa�`<�a�.Ռ�1�b�MLA�dOn��N�������P1sUuc�
׈Cc����\.�����w�.	P��*���[0<�n9WرciiZ��m���F�?$�m~�"5�u�f߹d��V"
��zw�,-��H�/�*
�Ů�Z> �>+D��E��󶢎�X�q�ݥ'%��$i���}J`�p!2�&��g-�N�g�E�C_9��8��Y��9뵈B��]'�^�O���%��8i�FǓ����ݢ�c��a�������)Y�/�l�N�N�h������r�+h^�촩j�=�8/ӌ����_f��-�޲Uh�R;�A�"�:��qU�}C�"�'0i�*���)�c��;3��0�J��%Ǡk:ˇ�_��M��Ds]�nz�?�;q3�ۧ�%ꏶ���T��'����I�cZD���=���Ӯ�!�`�E;�7k��x�	k�8bCʽ�9�/U��3[�Sky�Hݖ����5��l�4~l'z�u{>���yMZg�:���?�ޙ�K]��c���V��iZ�]& �|�-��i�̅��/$���i��7�&����H̆��`Rp� �fq��NC���S%!C.���k�2H��g�Fk�T����|Ϫ �ٔ6���}�&�px�N$:���m���<�[����i�`s��^*W�e�R����x����t)��~�K8���N#}S8�a.;f��J� ���
5����D:�+m]�M����j�U�vw�V�[�����6��.�� �����c�1+Մ��[�Z�3���Fރ��rߐGh����fbY!�B�����!��H�;D�0�z}���
%6��dtQ�X��2����Zx�����e�P#����6��>1,��q��b�u�O�)���i)|\�u�:;>1ϻ �i��@qcOʢ s~/r9D��ґ$�B@8!��FiT�`D���AF�ID��8q�R�o�F�Η�&�i�EZ��n}��V�%sI����$Dw��p$+��D��q�?(�z�S���*,��d�����
7�D����� p�{X�-]8�!�, xpke���;���_KLB���ݐ���mF���:����d��2��@�\���-�dlr�(�RY�2�5�cÑna��)���O�z_s��:T�Wb����?v�މ�ST�	n0�Ms	��mkO�7�5�?�W�b)V����C�~��Ā��|)Ԛh���K��O�L*]bT������6�k5M�����H��fv�����'�%;�A��P}�'�y���0H���	�<�0,����-Mp1�SV���#��{�'p<q?����%�Y�LK��2�=a����~��K��X������T�t�������Ѹ�M4||Џ��յ�X��`��ᗋop[�%\�� +eX���E{K3�w��1�o6Λpwg��.��2��C3�6�F7(Ul�>�9���㪌���tc\��H�
~��L̿"�)YZ�`��a�n_��G�����D��f�o�'�NF��1�Bp|�g�T8�$ǹ;

p�������@A�e���gªZ8�Pd��yt]�5�X���ٕ��3�,��n�g�,�A�/Rω�tY��/���Q�;UŢ.�.�nHX2V��%��{ؗ���I�)f���6f��-NEG�:��Jг�/�=�Z�&ͫ,��u�C2������F�g��m��L�N��(�_��UW��a��u���� IM@���
��Npj7�=Пx��������]��b���9�X*4r$��$���i�2��7D��B:��p��;�[e�x\�N�tt�m���}M�T��
e�g���ٶx䩶9�В� ��*���P�aZ�ŦQ��@&��������קcdXw�6!:��#��e���6� �0K�tQ�1k �'ᙺ��T���o�&�{� ���}(���^��R}��bZ�?#إ��b�0�C��M�l��ïk�F6:�nqO����������{Q���r���4�{�@*2�gWu�irQ���˞}UeN�>m�	��9 �㥑�+����U��	�¬b�P�gG7f��"��(�=Yti�Ro�����O%fiwv,������K�Hq�� Ϡ�F^�l�*7�	��'�-2QP;E�r�������yU9�o�%��]m���Fux~:6pDߢ:`��S��h�k�i�>W�J��ߒŗݻ�S~��G��կ���W?�;�LVp~~�LΡrh�V7P�;{2�%6���8TD5��4]�o|���ل�W�%��qP0Ű�:Tp���W��X��� ӯ����cW��V���:���Hc����%������RZ�Q���-A{�{�쓘EF��܄��m�23�
��*�����9k�a 4DF��R���1������J�!{K�;^�C�6�^6�C���O݌�����N�5��o��Z��Λ�)VE)�cb蟓mI��)���U"��=���k��B7Ok	��\�7ͩ/~	ǘ�AC
=a5��sB'W`2�|�/��/"���/�,vɾ�s��/���o���0?��Vw����.�A��w=�R,ك����a�N���^��IvP�0�Z6f%V�N�ۥՎ=�G�_]_�o��X�wS5n���!z���Eu�(��2��܀�qv�	=��ih�R�t��|g�P�~����� �Wl��j�nu�4�ʥ5*�/\ގ�k��C3�1'߁>=�Ib	�PTJ�;���G��"��+0��=D�`.����Q`�~��\�D~*;��֣
��-8�J�����!�-����)��2�HHP7������9��&�y��d��gɳ񒵒+Ց��K�z7��;�1�ƴ�������2W������S�`������uI����;?ͬ�Iw6y�"-��_��S��/j'X��]��_��b��O���j��ۃ��gP�..X���@F��
�t�ߔ��N#R������	XN���p"Q��qؕK&��ķh�^�N��{�Vq�X����g95��(������QP�ݷ�cj�%����j��;���<�;��ǒ��3�����r�m�P<�m�Q��L���I�]ǑQ(|�qr!���7��*��B�Lc��Q�����֙_{3���q3p��R�&B�5��y����m<�z�E~��jr��9^��f�&/Fe�h��~�\+mh{�Yۆ�Z��;�Aۻ�2_{;�E��!�V�q�y %�ҵ��ˑދ����6	���8�p�.sS����@X�N�mT�����@�Wɋ��j��U{j8���r�f2�F��\܃1��]�a�@�R��X�d�B�P�G�6�@;2<�0��6-">	)9��U�W�-0�ϐi!/�&��"��&4���(<�b����ro
TR�q����Γ!9|b��T��5_Q�"!X�,��R�p��]�i�B�����a���cX$E�UG����v2���m{��h�C�IvOͤ�o����;RΉ����:#�@g�ghcuɨ~w,�k#����k&���̬��/
� �2)1<���N���CJ�W<��w���LO�3�D�pjV�rpm�̰�ˌbd�K�B�ݖ�ѭǷث�`k$������4��o��R��.#���ۗ��,0���pE��J�;5܃}/��yq�.a��3H���$�R3�xuG�&��>,�"T��jd�Q4`�xl�r��Xj���?��]����}=�@�a٫Ա8۪�1ʘD�?�ƠtΟ!:=05�_�߭ʢ�-��2���=�G,o҂��F�Bb�L���1�v�1�Ej��(X|0���b#�wn��v�K�͘�������u�L\��\�%Y@�#�r�R�.��Y��+􉥭����
��M����Ϗ鱛�X�?��[���&Z� ����2($� �(��]u��J��.m�������J��F,2B�	Ù��L���7PS��K�D�va�� &Φ�}1F�L��u����&X'<��	��o�KE���-qKU^��f\�(*����
�uo�n=�ī�I�sĘI-�/ӈ�є��-�x9����!�/�y*�RiS��G �D1��ļ������T����F�|#�2/0�Rv��Mm�u�d�� ��?���]�ޙroź�+�%�F�1)p����r��
p� �*��o�xf飳p�����Ŷ��=X͜H�y�fr��t[#>�+>-3�*j����7|��T=�4z�Pi?��e��53�Zml`������E����"6r�'�)�fw� �h/�^A�};����.��~{dBLv1�v�ys�J�7�����o{BwJ�����*σ[G�n���*����Udܒ��E#>�Ɵ:Cj�v�D��=�j��L�l·{��\!��i�g�_ ���W�� ������hv!5<R�W���a"�
�!�.֋5t4J�}nT)Ւ�m�����y�>��FG�Y;����* KBLr:�Ѡf�؊���k�EO�BP��U���wS��=����ʔ�}�)z���	��G�����W	,�}"	�psÏ��݂M���� ��(4Y�V�3��M�\=�fZ�sg.���8#J��޾bRTSeb0(�3HT%`��-W\߱}�y&�$Y��������gkG�9Az2m�
��>b!�Vv��E��w�N")e����䟚�V��UI���
�N�'0�,�s��$� Ifz���jS��خj��Vld�� ֢���5{"Q���b�
mPJ,59�6�;��׍���ڗ1��\,�@^q��K��(�%چ.K,j��X�[�K�lܜ_!�{ObHw�; ˋ�>g_T%��;��"z��# A:Z��p��k��B0p�í�`��f<�I������Mt^M9���x�!x]����]|� }����4����C��QL�E(��jB��6$�R�N�d��3d�>���ޏ�bK7.��Tty\����&_����xF�g[�|��f�wX��Kw�/�@�V�����C�,ʸM���W^�^aj�Ss�mJ@'Xn�.ׇ֙jfDd�O�����l�vT�& WpQ��b�?Z��o�u�ދC(.�7!�{|�z�^�����gG�����4ɣ$�~��qdd�w�����-q���-emX��ql��eI��Xm��dq0R���*��X��s<�oɇp�!z�$. ��caz2C��l�ef�z":��#&�Z���䎤�N8�Q,93�rYv��\�(o�h����l��ؕ�t"�7��8�MEN��#��@g��X�ɵ,��x�w⌂��4�I�q�.�:+ru\<Pl�C�4��U�1)�q�>��i�1�`Q�
�NR~��FY��_��QFKg�����F�G��a\�S"�M� V�Ո�ܰQ8�z�f��]�{Y��D�����K��(p��HA�~��R��I"��hQ��� �փ�f����PJ޶�&��l����o�(y# 7���>u���%6+����?�G9�F��1�6b�W�3�"�N��6��Hٕw@�AH^SD��G'���É�Q����'�vā�o� �`��ug����*@2�A2Ӂ�iϽ�oy�)F^8���[�w�\�m��]et���h�1'�n$�r :��To�1s#�8;�GMBU�(MO����}qF �\���\܈7"�%e��j;q%���l�?b�[�M%��Isr~�7g�3ya�_ᓮ�0V��x:�9Ҥ�{fo<�KQI��A�NJ��.ph���8��	1Am��w��8�]�k7���2�����:C���b��D���,��P�uY)
�>Q�=�׮���t�M&��4inSTzg����}j��F?��d���cL�Z�|�'D���܍s��IYNC���6޹Qs���ț�=�x?�'���`��e�b�	��7[e�=/d���'Y�����$l9:��̤��{�pT��� \�@��%�?�z^n��>�_�cx�
u�B8Li�z��P'�=�N|�
�2�.$d�H[�
�� 3�p�-�u�-�XTҼR�>a�n&�0�)��Of!�oA�& �O��g����<�]���]q��q�$�&X��Ė4xFf�(�tgz��ʆ��(������F��}������3��'m�N-��d��qy����MH�^wYr�F�����ۼ�{�U�
����������)Y߷@T<H��J4�*2	z�V����l�}�S��c��ax��'"�Է��h�����MY�G�F|�q��Q@UtT[,6�/UP*�^E�8�)�� �H&1TP���R�A�R9��[T�րVa�d>��L��9�6���=�p޾I��/s�r��7�IT��*��)Ͳ�x �`�r��)T��:(א3%7t�2�ϕ�[�t\�I]�4���Gpt}d�UR��l{bn��D�c�.>ڨ	�����B�*��jՀ�����'�,���%�pk����`��X�Am�S1�o�n���#���!f]1�u\<�ق������c�b�����{+L*$�-�H\�I�����������ނM��'��,W.]���ߘT�#���,�N�Q1%]���6�j ��5(a���e��V���9*׎aVa�x�����m���V�N7��F��D:klߢ]��Cg����?�ڡg1#C��+չ� 0ℷh�>�M�C��b�g�'zt�hV�;�ɾ01�˯n٦��ɽ�-0����������_!�����f������iq���ޅ�0�����ufz���K�*L�!+�2Qf�5Fh�� nMj��L��a���׍���� N�)b�Ѓc���j���r$H10��������	����i�V����l��������:��V	�J�yVq�?�\h�L
�g�lw?6�0p�5�U��|*����EȍW(ԵK���<���� /�f��H�Y�: �6j$"�G�5�"�p}�	����  s/&ߤ�-X��x)�T��/��ؿb�ߖ�?1���g�KgQ�IY�;��Q�g":?<L��Ӕ�
�#�A���sS�p�0�L�����?����9S���;�$T3�b|���K�Nƭ&�����M�b�ҁ��8��W������y�#��>���e���HZaP֬���^� ���%m�[�t�WRaW�2�Oˆ��/Q�������D�(�<,{!R� ��"�Bm%9��ޤ A�t
J��D�|�y������3k��C�?ʏ<`�7���T|��´Ȓ�����S��%��4'�� �SE2��X��czHr2���1�|�r^R��]��{t;LH<q0�罘 ���٣��`AJ�]����wW��}w�T�D!��.��&�Â���#�?L|�,q<pP�_h�4��E�.W!O�5������蠩����iY_���7�z)h��4#����?�*�E�ڵ�<�zt�����10��a*�R��������Jf�a��S�\1k cg�g�E�'x��^�}6�~m�9������u����Ǖ?3'������54xay\�*b��Y:J�z������"�;�:�CK��uD�!-z�NC5�Ɛ#B���ܓ�?;��;&m�� �'��;γ-����s&�u���3k�g+��U�Z��_8��1Fa�K��0ڔ����`���U���c8DGg����-��%=��.Ga�S3~W��Y�r1�܇���Uֽ��ec~f�i��������nNUb�;�_60m�=�dsw�z%|l��U՛<��'��0��OD��l�S��1���:e� �B_D��E����O���S<V��G2{� b6y8�,�z�0hV� %�Y"f�"��$젆<�jS���r��J�V8�[��'���a��.}m,F�sG5Lg�(NZ-N�	쩷�5�`3��3��@2��$L�U�0�~+��ջ��;DHF6�o���GA�ܭ���me�JZ��?<oő؎U��v^���3!�GS���"M�J��@�ǌd.�_������N���`w���8P��vĖ`��T�>�Y�R�l�6b�{	Aƽ��}���f�%��o4-�ۗ��T�lx���o-���KW�<�����ƌ�2c��&fR��x8u�h!/�Bz�� �~�yaf�g"�
�=�s?��]j�J�u.�E��?�mvn�ʺ{$����&Y=<r�3��@F��ڋ_�$��ur?ﯘ0�R�v��S�`A�O����A�����@�L^Jq8<�F*��3<�]P  h4�~f�������@<�9�@�#�d}��>q�������/c	~$��RG�~nk �8��)_W��7�j`Y���E�i� E��}�� ��R�E$�m�җz�^�
��(J��� %m��S�6��I���J%�8,�J�n�*���ج�7��]&ā��QQ���AIG{.��-�a���Ȼ����w�`V�-M�<�R�V����|t�j�n?I�aI�6��ɦM`�	l*bUm�{�8��=�J�m"@K�������^�J�a��*K���R�W�PF�P����1�#s����Gn�ݱ�`'��������v�#}uFN3l)��qWF��[�0�$�p�K>�=�,�{� 辌���_��R"��I(�)��%<�����wz�R\��=���W��L�m�����d����J�0� � �_�G�/q}�b��&�DYkAi��ja��挣��P�\ܒ=:�%A|�2"�eZ�����OKܵK
��|���Xu��<u3:�.Q0'V�qʝ!��z�����>L��TU���!��A���7'i�a5 H\�	��,Y�S)^6ޓ��	�ah����2����?ߖ/�i��!
"@(�S��n�rl��RQ"�j�,K�KFf��(Ǭ�$S��]��A�m�x�Ӭ!���  
8��,�R(��ֆS���eM҉����7��{Gs��M8~�l���Ĝ°0(c�����OW�@=��s�s�ec�OmD]�����k�E���O?D�t�$�҉�s&TW���)R�Hm l�9�5��w��?�]�߾���~��z%]II��N��d����E���yLl��D�L7b��M͏F�P�ҝ2c��[��6��-����)�*�`R����w-{E[�R�hd���s�4�r;�����s]̕����{��$�{��:�[اjM&���q��5���%�d��!CDk`ږ
���t��0N<bB�ۺ۠LhN�,9��sO�0Z�\%O����?��B��w��l�y� w�>E"�$o6�.V�ԙ�Ms�V�ɰR��3
�<�2J�8]�$��` �s��v#Ç�oT�
l	Ձbm���Q��8&y"�G���<��K�T�糼	p2N��*�:�}�0���u��wW<Y3�A�V?Ա�������)��S��C�D̄
"}�I0�Vu��z�Կ���h�|�kw�w3�Z��ῆcK���!0K�?r.��[��EM�'Cb)�/H#���FAt6��e�S������
��i?�z��-�o����\���xD$�&�I;�,lCǘ����P����K-db���Y�����ҕR���y3��Cl����Y؇�%5�s�:��S��beM��5ı�-#�=%�(!��;�<�^�Ojc�3�>�]Z��:��D��v�RZ�Z�h��O�9��q`4����/��%󪐀V�����Ѯxd��J�	6/��
��� 	n1���iAT`RqĭA����56�A�<�z�$s����v�藛Sh��h�@�F�b�s�;���-��F�	a1�"9�&h�^;F�}�ycUq.�*	a9~�Ldt��2�Z��J*�m�y�X�aB���;xU,�L��J?�zn�"���Эp�@p\�wK�o�t�i6]��SV��v�-���h~
�Z���!	1��`^�\)7����3��\Z�X�4 ����=��6t��c����&� ���+o?ą}��{_FUϹ���_�s}Pe���ӓ8������͜
J�R�RXr�S�6��~m�ˬ��<E�o�)�0WQ�8ja*�gHt�Qc^'%½�,;P�L�g*��.�6��M�8����
TO�GV��K7�+tm0���+2�olF�rh]�T��XD�Wyw���}~�b�-Q�;M%wv�@��;m�V93д�W$E$S����^T�z�^~�E��~v,�0�rR���������W������o����Q�N�����Yެg�84P�y1�1�<�)��B8�sAw�d�q�kg�J��k��x!�PI w�3Kۿ΁������s����r�b��׮|=��r�
-%_�`��%�ס|
�31l(�� �/��Zv��3�*����󩞍ulvB�Ê	�.���y=Y0��d�d��oa�*vjb��y+k�k �R%���i��ޥ|�]�-,n�S��pg���Q�ʍm�Ei?,|�6��nC����=/�sc�iW�W�Tcd١��Bho��Q
|��̾�@��B�!��xA���9�h��|9$�rؚOv�*�I�i�Gܟ���ҳG���E��2P^�1����LY��w�:�ƧD�#�>Pl&cr ��N��#ޭ�Gصdq5K���%�)���&����&N��D��hSvEs}���; �WE�B�B� ��# FBnY@�z{��I��w<]�ח.d���ITj��~&���P�\XO��m���)	f�#I�A`�1�^��r-o��uP��c���\-:ݱi|R�7�R�,������;�'���g|V|~^�~sO�Mu�*�����ˆ�?xI��Nxĳ#u<>�Q�~#P�a�q�@�z��;>e�&'���c�-��)��gu��h��(�ܤl��\����d��O6�b�����·H�׌��~"��.C�@������:ڟ���;�U7$霥B�2P�J@�d�ԭ8\���5�}R��@a�o�DH�$�9�{��B4�����ri�)�������ը����ʞݻ�$Pv�Q��A��Ȥ����l�_����`����f��G��P$��cU�p���n��5E�p�%�	� h��x�o�dC̓:�O�s�h%��H�6�%���<+z_.%s"�c�L0��,��Po|_���p�*� ���W�~��ץ�mF��t3h���f6���6����L���aپ���J��'0:wb�oWZ��Z��^�P�_s֜�仮�*�#ƒH�_Ǯ���JW������.Un�=$?8j��#��#)߁�Y�9����
]'��/�Y��{�L�:Ӌ���${�G�������^��.X���f��i:\�����x��Z��