��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���l��o[��ɴ����>�$��	6������b@�	������b��VJ�o.y����L4���Z��1룠������	�<�~���E`��-�R`��k��-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_d
�t!���N�S��گ/�TNM{�C�5���M��;����L�S�:�{���\p<��)�0W��B�R<Qt��Ԁj,3Ӂ�v��`s�HW��眣�U�Z.͓k����W�z�N��VXi^�p�ޒ�}�@\�-1���:��[�e�,t�^f�>�Q����ԍ��H�Ѹ�C��!K�1^��C2�5�V
=Ҡ�JزEIStH�-��B]�2��zs��yt�I8����J���'��z;m�\�{�����̀��N6���@7Q ��>����@��E��
f[l
&e���9��`��-�m�a�Czq0i%�;��A3��U�Wվ�f~�I_��[ӕ���lT?W���;��>��^#N��D���P"h� ��2Ӥ�ĭ����Y�5b�8\�D�5o-Ƌ4mX?����J���8	+KѺ��M�U9">wi���?[�ͮ���9��k�e�Z2#r��B��t�6�����j���|i��W�F�1��zG��W���yȂt?�۬ާ��CGS��+�
.t�nP�0�]�t��Κ�1�MOx8�Ml��v���6b��
�S��2����z�]��L:F�켭�p���
�kݰ��$�ِ]����ma*�F(���?���FFN�t�s����<e��� S(�jqʐ��QQ���_iz^�̨�)�n�?K �vv�b���D��d(�Ѝ�%�4e�o�F���%δ�����V)i���e������e�I��Q@J'��#ؘ�&/D���j�~�y],��[U=��I���}���K\Zd��һ,�%H���,�d��G� М�q�u��<n��X�D���;���nv=��h��s�I3Cs�ti�ɰ1���ϻ�g���mJ��I�������]�,0��
���_�]e!��R��Ouy4��	����T�HL�Pa�>9�]��2��>;$�{&�EAy]��p��wR.�U��M����x�xQ����*aV��c��rD]�5X@�����6vy���R5���Wi�M�?�?��@�-<Oވ��|7���ce%�팘)R���S�$p"���<8����G�	m�ծ�3�<C�m�"�&�<ܻ��[����E�NKlh#mSg����<kt:�*���o,ۈUg u�
�ev�7ɓ�����:� Ԟ��m��\GX�[Ձ�/=���cu=����8&�)9���x��Zn�v*�v����S`� Ȟo�Ť�C>�җ�v4\��{%`�˲`����.X"e�@�f�wx�����|�݁V�$�{���@�#5���:Z�nja�B����A��L���`��������*��b�;�'���.NDZn�P�j`Ys�<���E��<:�<�@µ
��l�a����Px���t�:���>������0�<���������� �������Ej�|�	�]N �][,�4�Y�6d�
��&c��T�aLҟ�鶾��r��#}�i$�N7F��g�h��"��D�;8z1Uu3JW���Ae����������,^�L�+! ��	��%?�A�y����f&|>jvQ_eN�/�H�����h�;׸�os2sW�*�%�����/�i�����'{5��*��]*W�UY1Zb���7O����~Ԣ)]�O�?��.�~i���{�+�����#7����r��c����C��vn�h�q�}S\V��i�ow�J�?|�[�u��sg�Zk�v���"�쯠��2��4�8��&ba߂���7ۻĕq��#9:dEFe�Q���c=����a��g�haɶ%Jد�5>��ݦ9��e=�.�K�_�Z�Xd����Q𜥛���P�.qķB��P��-���8{�WR*y����
�Mh�py�W�iǶJ>'!�M񌿢��99�X{���F�h/�$"���%��Z�Z͛��r�͜7dO������`]�漶�X���'�'���y'�fΆ��[&
���Pu�7�b�*��jy�Vd)�����.c��x�������L�l�,�Y�NA�=�%2���FUJ0"E~(%C����H������/�`���&6.���W�&C�%� khX�ɖQ�
�_|ԥ�����{�$�k��Z٩�3`,�]��QԌ��;�*R^�tV�W����rr���QE,�,"e=��������e�����<�7v��Y좕�"��د(�\]\�ŗ��]s�F��,�݄�ۺ<��,7O�Znc��g�U3��� �,H����pte?�'�6��}�~4���4�m9\��"0����K5e�F�S���W�S��E�	���V���@6,�Ka�0���͗�2G�$�� ��4�1����A�OHJ�}���|p�
8���xXs��\DE�ɭ��G��^j5���Y;i�K.3?:}�U��ㄉ��p
g��7O�z1�l�A7�� �,�-8DG�4���3�������2z����	5K���5�yh�F%�MN~�]��@cY��	6,��6I�g�M䃘��vvJ���۠ɺ�fA�����(��X�����u�f�|&��l6X4������t����`Z���OZ@`l�]i�z�����@�8�� ���N�e�R�K3��<�a�V���O�����Y���v�ze�f�������������<�, ��x ���_�$)���W	�Z��u���x^n�8E�K<붷ͣ�%���	GX�l3tg����r����s��gX0�h/��{�-�!t	;�%�q5qL}�9�7)X!0����Y#~��$�y���^y�c�P#���O���\�ʢ{��+'��b���詆��d��[,��y��p��dgu4�H!��,���E�*ۃʍ4�u��;&�Pd+:G�i�"7���n�^X�u2՗X��m>M�R�&ޛ�w�>/��vA�l��?Q.�n|�����f�)^e
���?�#��?<���!�9�TGE.P`��0{��*-]b[�l�tg�J�,l���i9_z�X�oy���%��r	l�vj|rsQ��+��s	�_��0�\l���M�ެ��F"��Cr�q�$����H�ռ�eS��T�ǱD9DЀ��x̽3�)���O��wǛ��9�I�\��=�U������+��;p��������A�dZ�������fG�1�"��ĕ"�s�V��Rj���7Q#�RK^Н�v�i���l!��B7��F��aʯU�3���z���Զ�Z��0T���[�ZԚ��w^�g�Ȟ�!�Թ��B�\Gf+�	�x*�'��P�6�2�ƠZQ�W�C~"��Er/���Oձq� ��Y"��|�����v�]��)�+�+�>��/G�	s�p�	;��[�3���<�������B2��}��3�W�Q�A��� oCny�^�E+�[�pTP"�̙�d�Y��x(���C��8�/*��e���%���-kz�4Pk�f���*p-0*�Y��^��n���v���vY4�ї���]k��3��Jn�f���ȸ�H��4���6�g��wQ�9�i���:ܞ�;7���^��'~p5�Ma<!�||Iլq J����wx_��x�){-n}I���s0Ut>
��Xڒ����6J�P��^\�����v�c~��8��%�1������o!$�X!6�'(H�����+��z���Ni�r��3�����wT&<E=�
�;7�h�^�E���3p��nؿf�ry���O���B�h������Z�~�ߒ��6�"�c3�� 8�:��s�<�iY7�V��W �.Moi0�ǳ���}���m~�~g�w��~�)����}��P�}��p?z�r��'�5������0v�_�#�<�^}�Nqd�իP�Z㒯���CH"�\������=���(Tl;�93O�ߡܧ)�h�g�e��0�8c-�="�Z�E�V��s�_�r|f �DHJ��"�<��8ו���|�Y���f�g�Ӽ�{�v�K�~���֑����SP��zt�[�	��ù>*���{o_��!��{�-�}7-3"а>���O�{�T�>oMJ�*%੦��E���X��1j�ҭ�k��&Į0�{��P��	j�H�1�K�E2x�G����E�݃F�X��#�T�	@��'��v��h|vT��E!_��F+F��"��̘#'J|A�S9�iho�g�2���7?}��DG��4o��3蘞%R|^I�{ғ��{��T��yJ�f[��o�e�'���������Ԕ�>ky6��D�7�3mgf���(����6RI�
� �vk4d�(?�r�yp�r��4�9��y����b�I�!�ZNA�B�LV����"*�������t��䀱��V���̲w�ܹB"�#�*��1�~�G����u��9���N!�_s7����{Y���8>�x⎍�e=t�/(�r��G������A�~|J�}K�r�΁�y��1Y@�P�_�l���~���e�4��`��B����c$�h���.$4-9z��G�94�o�M�?�&~����8�1+ӧ鑋�ae�,f�����nf������P��,�6��SD�UK
_V��װH$�\<@�y	v�@Tt��
�$V�u&BNA����n�XG�<*���T�����{lj������u��ߴ2�"Q�����0��P�����<m�;6����0�g7dh��!�$�Jhʋ�'�����J��A���Rro�J�k�ѧ��%�L:���t�I0�|{:0DX*��V��N�\� r��� ,��|���{��.�5�p���{��Z�)�Qu�u���o*t'�[{�Uܞ���uҮR4զ?��چ�^�].a�jW������2�jb� �j��=t�V���Ճ����K�,B@dW�ײ9[��SEݭ��/�������'�O�Kn�dU8"I�)��o���Qu��Uۡ-[� *�ۿrbq�O���L�W��} �^��4�{�A�ܓ�S���f�j���)���U�	�s��!X����ʻl���L��хF��g��,Iag�V�4����*��$O�Q�Fjox�Ք��Ft��7y��C�C$��p�-���Չң���Ӎ��)R�q�DN�z�(�����<�7�7��s�D�;��j"_a�l�j3Y�NҖ?y���>ٺ	�*��\�Ĕ�1p8�6�{[4��E�;nKT�`_�@{��|����J3۟��@9/j�_غ�u���eGP��,����\��5��׸v��LIe��B[g]�S�tT�����Zk��W�eU�vvzy��E82��F��P�Ւ\���I1�f���Q�yF�����v�Gd���u��pʻ����� Z �ܡ��[2#ń�l��x�Pv
�f��k���w�����b8� z�bT���f<�C�M���N���sS�ZR s4���6T-�-֢`BN�ɵ��$t`�`emv���t@m����֨�j��\=���pȞx�/m��Fm�Y#�UY�	��c�哝u��������+s`/��4��M�[A,,�P~we�,>,p��f��>1�=��� �rcq@�h[{/~)�p Nܯ��W�y~���"�4Y�"a�+S�0X��2"�9��ߥ
���r=6�e�Z��	���v��,l���ۑe3I� �!���1����^�����4[6���H7lP���0�Fն���vC$��1˻A ��1h\F��O��_�jxz`:���ƀ��N������+翥9�n�����K�T��d%6����R���j�-���du��AbL����D�TL�����2�.^��rd4�1v�İ�I@��:2!\"�!]_�;2`��U�^;5�`C��*"�e)#IT�Ҳ\s\�p��g1��OɇZ����|��z�u��5��{��3�r�.�qQ��z$i�8�w	�����P�}؛cI�tu��m�����!Q_U�r~:�z���}�h��.�A.�_�b�o"N��l\ǎU=��և�a&�́�}e�<��F�H`6�~� ��k`e���o��,�wu:�qA��`�IRm�'w�e��v �nX����N�QF2�k�\��YA׷�p����J��Ec1�W%xu��rR8l2�fZ��KjfO��@�Y�xF����+�q���.�!�iחZ���(O7|n 1E�.0H�v���=����u�4|z(k�T��T��V��G��Z��A}EJ�����������^Y�f�#2��(C8a,=R���;��DxZO� �З�z�eW�U�)6N��,���?U�Y����*�N^a��?��a�WdJoW����(����B�0��s�v���a��L 5i|(w����}�^����֧���9�����4��s\4ir���vF��Ԃvd�iD�� ��B�;�D��b�O�&c�ev��f��ɳp�yz�t�d}�^O���nK��@�n}�=�w��\��L��M�FJ����w\i�Ǿ�/��o�7P��ũ�i:xK~j�3��#�;g��ad��K>(�2�-�uH�0#����r5�,���E��7�|��Ϟ9�M���P����Ԑr�5k%��ݖt����\��*fM�R$64��}�*۰-�P�!�z�#�<K ���I��:;�ұ�/�;Uk�b>�ɪr-p2�v����R{a5�e�? �J���<��"g]ǃ8 �U��a�2�	7�B�۫k��:on"n�,�����)l�B�h�_��>��9�)�5!#3W!���;1�kȤ�YL�5�F�^�noNv��N2RZ�Z�t��C�6~�W�[�̄���숹���Ŕގ�1���0��aF��Kb�n�	/
[v��Ǡ}N��PU��
�a�c�ra��7����eu=�*tȾЍ��3?�q}-lwAF����3�W/?����S	��/�����qor$��	*�vr���9mWt!6DO��$.� ��WO���O��5��gH�ã���OT?b��r�ټ*u'$6$�Ba\ڷE��Ƴ$���~rmZJ+8F3����&dS��q<m	�.�(���1��W�,��/s�:'*:��٘�]�����5]p���L�s�~G7��ZC�����-��lꆿ�ܼj�Eh*d�L"�4��1t��>I�&�]S�s(���*t
����Q�J���-A:�ؐ��n'����}���9M���#�8�n�f"�qMo�A��_��8ߞ�Eg� ��O�Xa�!���_��?�5�X���U���zȢ,�*P7u� H��f$8����-��ð�O�0�$��z�����=J�SjA�0�H�8F!R��'w�:�ka3�;�����JY��y���Ӄ���	r��8������yԣ�.z`8��s-`�Nu������S�R��9�I�H�&=�����p�`�!v��2����|��â\V�c������|{�M�>�DE�j�o��趿]2����&ގ���U�?����Kg?��F��6
~k�~7�<f�c{���ڧt�a�Q�;`�iDZ���,_�Voy��8@D��u��3d�������Pa,͛��ś	������Wt���.&�A��O��CNU�am3,��-�XLl��uy`f�3�A\�+ƒK���ϝ�boS��0k��v�0��3e"�A��W_��&�;Ke��ԃ<��bn�w����54\-�@�7w]9[q'LZK�_�^�v�"�������7X\l��]Jk,3�fP<]���1î�@P2�l�>�D4u�-&�����x�{�B��r�Z1wת�*��3��z2��(�u��׳wJ�i2p=��i]o%���~�A�M0�k�d��BMvV�ni�>�&�莗����W�z�$<`�`~�S�}|�a�����#R�M�d�g�]A���m����o�;���`�Hs�X�B��0�]m�*��JEM7�\�./�l��ϪmlY6�&�I@Zn~���m ;���	M�*�X�B��YT�O}z�������5���-��,��II�৿H��������`�T>?�{_���8ubW���;���:Q�da+~M�&8�	�Str�y;~��q/���9����\���fiб�c˅ѝ�k����~VM��6��K����\���¼�	�P�qP��=�x�Q���ݟ�@� Ǯ�.0}��ٲ�Zbg���)sY�@�qx���
�#�	��;^�T*���]�J�ԋ�h��/?uː����%Y�V�j�]e���v�M�r� v3�˔���W|�F���$�Y/𜇪/��^en�.�͸�G u!�[��VK����R:����W���m����a�f���§i� ���]=F��C��C������!hu���2��or��5�ts������ C��r,�Cm�!H��Y|���u�D�)�+\c���(��.]��U�0����K��B.�㓺"����@���D�$����+��>y�S��d�ݔ�@��2��k(�02S����B����ւ=�]{�)�E��G��|0$㇧Hg����%��
��`y���y=4�o���$�����tJ"A�3���I��4��¿���z�Wsl̻�CQ�T�v4��E�*�⣐+�݃)6��;��έ��h#a��_
f9Bh`�2�9	���,K�H��E3'�j˙���I���y�{�n=gsKf���k+U�-���QDci�1�^o=
h�|;!�RGAiy��6qZ��:�-�%���Ρ���;�տ��-�u�7�\���r0��~$I�����Y������Y:�ݷ���Jl.�ɅF�tA��j���[,��� ��`��P �:IbTM�	�� ����g4ʖH�lŠ�ͨ��Pe�@�$�Y����|��������	��ڒ��krhD�����&�0T��,�m�w�TU5'�b��L7��إ��̔��7T��
}��T�X��[�x��ӯ���l"�a1��nvcn\!Eq����J�|F��F�B��9�i�Y"�J�_S���fH�ϫ��K\�V��G5���<2�;�l׳;L�<o$������mx_�7FS��r����L�?������P]�;}����uL�p�٥�2��&��ԡ�b}� 6M����6ޘ ��\=+���������?"��(�p'5\u��E��I���MT�f|����{����9�!�W�3W���+��#(1R�+�~� �T�{\���Omԇ�JXfWD����W\����#OnpM��X��;P��<��	��33C2u���z|�D'�ܓ��28��sƬK��h��i�(OSZ��po1��3Ni����«MKxZ��uD�u.P�)��hG/8N�v�^h�K����s�m��o��|�����-���6� })�W;;���yg��E K������^C�?&w�j0�&&�����hձ�x赋�J)ׁ2AC�x6�<�Y��B��}h.��e�~�@&
u����������u��ü�$�W[���C�).�i%�v��YWy�^�����mk��s�"�A��z����	O�� �l��"��:��C�_����(�cٿ�����j�l��4���u��uU���}�z(��$�|����:����Li%�U��>�:~�ȯ����
�"��6t�9E��`��EA�~�^ʥs1�q��k��;}��v�5�B�G%���N�N��0HXrf_WR*�@�_����
��O��$��漤3�{���p�>11��D'Qq
��,�k�	>�B�/�DG��2�Ɠ���� $�q��QtX����32�����U��%���Y���#�=�K����^g8�U���GO襅��tੋ[��qK�:�ф��8��qA��?���s���m�)�Sʏ\�,�
���b �m��m�/��z2=�N?���z5��JI5�'AOÒ6� �h_����-�ZA��� �nP��&����}��1v���W���2�`�$�3a�wv�0�sLc'������.�r|<Q� i����(���X�?a���Ԡo�\��6航��|U;�F��MLW��~TV_�W̶��Z�
ʏصM�p�+�;��ۂ�ߢY�j"_؉3v�xų�Zf����������$Z��o��n]���Fr��[�f�\gW���I��v�2-��WG�6�'�c$��+j�@3�rz�g�6�GR<5�ଣ���^�ς�/vR��[�`���ݘ�����5��@`v$�aQ*�����3�_���($�|�����v�o��հ9���G��~��Y�O����c�lo��ȼ��JF^�I�N�J�0�J��L��k�(
G���^�H9*>,����od`~e��&4��x"�vA^�4�_>����^<�Vq��%�q���} ����E_�x6�h�tޑ����h���:!�+-Rph���&��\�!�ӆl2���.E�\���u�
C������l�y!��ǁd0�E�~��W�F�������{:6���?�.�L|�Y�`�ʙY� {�uȾ�c�5"�2�Ѩb<�jGL��9�0�

tλ����;ox1��h����X^ҁ�C"Cpð/��8m�U}�o�m�j2:�?$@�ㆰL7ӫ�Po��/L&PΥ�q`��a��s��O�,!�7u�<����2��b\����H�U���A�m�\p�@`
�`q�Ţ�%!J�ɰ&��#lh�rj17�	�6gB���ϗ�ApJ���p��)�[�X�xN����̤�I�{�2����tߤ��<:�og�"/qsJ����ȝ!k�\�f����[4��~9�t�����Y޳��.̽2z�Ҕ�`b}7�&�����z��F��p��&e)����D��1��Jm��4xס*l�y����<J�3�x�N6��@Z����U��#�|����i��~�n�F4��ɞ���z�K����a��ӓ�S���k|��0Rλ�����I��]_7L�b/�y㐼 ��<��Mj��2Ϟ��/ڙ`��&���4���	e֍n����Q0�0fy�;3�"x�1b{�'�+}q&�ik��ͨ���
�Z)�Y�m)���ӏb�'�nL"4��������NSwf��Ҥ���s^�t�耺#W`��<@6��Wh�����7�d�I"�8����f�Bx̲5�Dl캭6�+�����t2گ�?�f���%x�rD�4{���?�ټ��N�.��X��� �K�s6�8�0'>���h�A�����s�6��T?��SQ���y>��ϛ.��nԞ8�cGyS_ݔ��V��M����x�Zޮ�(ߕK�@��x��pۊ��Q���l�b�(Plf���T�sKa%j��Q�q���]?%�G�L���(��e*Kɷ�cO�@5\|@��o�{���d`���GR�����:��ɶ-��v���&���sԛX����4�[��a�t.�C���m9_�E�m�����@#�iVx���E��)������i��ۢ
un�;�w�֣����^$�R�u�R�AL�l{
���a��;.��PcW�6���ga�R!���P8ɫ��P��Jk~���3a��-�_���<�p���/�?Ne�c����Bk�o1	W�i){xyǙ���&��%=ښ�[�
���/�:y�"h�0���$����P�t�א�;ڳ��AkF��Μx1-&�;��`�x���F�	A`9�p%����l�0�O���`�W�Wt��v�;�^����( ��rOb���������ThH(\(��0�����h�0�����ע�p��\Y;PX�|Z�����a�����{�2��)p�v���l$_/�"���o�1������C@G���� �[I�W4R��Tۆp����|ܢ~'�.g�㇥/C�c�&��S</[_���]+4F�OP�@�rOZT�LP��h�#���+ ���v/��U�9�~�*����Q&�%.�N�~B#�{f���{�+�|���ed�B�i�
 �T,t�D7�<�q�����`IsH�����?��N<A������1�їe�u�s�[�.؃���<�r�	��#�mp��N/t�_Y�܅ƀˣ	5��2�&7&��Ǟk��<ڽs�f������뿉4��t��q�j��i�Q)�+��e�i��>7�1�;��ҳ���;i	#Oq�l�8i1sr]93�B��v�L���(�Ճe(�o�
�P����Ɣ����>�7cXʖ����#��!�?ۀ�O>0�V����Q ���i|���5��s�p��l���-\����r��v?�^���c��H��T�w�BMi� |#Tòn�	P�A���k^� z��q�;�)OX�Z��S��D�"�]$��2B����?Y�� &����3>�[^�� �ŗƵ���uI4Pk�83K��W{fY8֖��Ht��ҍ� ��L�kB �x����<3(��ĉNd#?\i��[(����>��ơ�MSjQ� �ϊ�֮�p�kEi&!J�4�/+�JO�Beɻ���E0K/PJI��	�`���/1:@Q9ҕ������v�,F�$K�H��\���	gB���P̘�Q��Ė`��x�+���C��K92�� t8������uJ�=��ZY�Բf }��"��ן"�|����ӠZ��R�4�W`�s��A07P�3�m��88�ǑZ����M.޻��BN�[������X�б�	,�7A��h5j���8s�"�!� ������s�� �F���)SX(�ܧ�?�a@B8��f:0���i���5�,^��嫷|�T��ܨ��0�B���?��w����c��t"������ �������ў1�R���GH�m�K!h����G&$s�I(M宼ۨU���ӓ'�h��+ƻd���.g�:������u'?�q�ٻ����m�*�C�Km^֠���]�^-�ܣ;��L.�"�T��"p��%�M���q��[Wp�SBޱD�;!E�G͕d��{�T���>�1�@�{3m�Γ�}��=�M��U�#M�#�63���1Qm�盵�~Y��u��\R����Ʌ҃��J�z��3�b쓤6�X���_�,2P�\5`0�Y�7�Xo.Nt��d
�9a1ܭ �A�U�7��d�o!ʚ������v2���%��5UH"Aۀv�k��n67;�`2u���j{�h��^z���hv2?��P�S��+�| u�`-���k/C�e8�:�G0��  �s)^����r�����*�!�W���#ys+�2%Ɂ��z���zO|
�|��U��V�-�ZE��W���Y��� ���cѹ���Q��/f�@94R�5�0/ �#�f�0`^忋�Д*��k
 ��d�=�G��'��hB�Hk�b����i��%A0�����0�{� ����u3y��|��\#+0���%��ڨ��9�f�{��+#A���n�~��]�8cs'�S9CU]
m r+���-�Y�g��p�u'q��R��qO �07�x�dj��PşY]]�ܨ�޶��`_Zm���S`��1�?b�ea&�V�y���Q���k�7��Q�=�a@M�cV�p�	�7�-c�W@9�X����60$����L�#y2��V	�������m���[��=�`%��:�1žT8�_��z��CChN���~Q�JՎ�l=�sgW�X���3��.���^�gzY T�z�w���bv��J!њ-m�~��x�v�5�R.n��ޗ��ȾDWd�Jg�\j�9?�PȅH�mJ�(�����W�ީ�[���D��b5�ܬj/�Bp�q։�j~��>���6�u�GQ.���u�^���gJ�-D}�ou[{,_�ν�ӓ��X�py]�J�@���'�;��J��9�@#G�W�V��؎$ʆ�NT��"�#��%�I�`>��fX�A�e���r����4N����eH&�F��Y.����;�af�ST[Fz;�Y��G����jؿP��&>vt'�GG*^����g��P{r�ܫ�8R<���\I�"0�F!V���t��Z�p������j�ѽ��>1��J�1��?��76z��kǥ�Y�Z=q,�-��3+I�ǸX; \D��lNDD�0��Ӆǥ_2�
X�����)���l.A/�r���jBA�rL"p���͙TIT��z �nE�����Q���##ԳF"pm~���B�k.�0��e��y���G�N�Z��"�Ԁ�΁����Sx�B���Z"����h|��[+�����B!�� ��gaү��9٢Us��A�!iI���R�*sA֕J�!�N�'�H�^�9��M�!�]�F�P�E4kUbQPIXCA{J�,�4�(�/�n=j��oyU�R>�@6�V���<&��,Վ�g����]�ս`3n��� i1�m��Zd#�p�W=`� ��dX�U��;�{l>�:vN3��>��h��4K�nB��pg:I|����4�����q	a~���,����w�]��h�v�fF*�\@d-Q�+ey׹N�1ŉ?ʋf3�����#:��'�m�İ�P_�Ǳl7��Y�c��-�=ﹻ������Dz���D���C��'z�c��vS���p��-�D)b�;��Km����|�@h)oŏm
��f]8�ʥ��"�S6����Xc{���;�O'��<�&�{����D���"Y�Cze �^esLq),����! ����Md���,�&�X�v��e�S�uR�&P�b~���ɠ�e��:-At�2�)�!Hɒ8������,7���E�g�J�C�*�iQ4]��O��:ٸ����P�H��|�$�a�j��b�������^xE}6�A6�ࢨ�Z4�����*�I=88و�w�HV�7�����f�c�J��ˑ!K|�$�{���u�k!�2Qdy�:�E͵6��N%�M߉�<�B�T��;}qL?Eep��X�Aj�k���r�	���P��9E}n-2[�����.�4��@V
e�DZM���ˉ�B}�,�t�-b�o;���"��k%��i!������#����������f"��?���FV�
���x��k ���8���˛�D$r������[S��������5�83�`�3z�D�1�K����U���+7�9]rtt>Y*o$&��gb����F
O,����֖���$�<1�o��Ix]�;-�\�oݱ.u�[͵#��G3��a�q�#74<_�4`�C�S~$�	]T��������n�L��|PQ��tdV�&����`�\b�q��[&M�`	m�<4��b���5�Ek�j��YO�v�j�]
:��y=��SnA��ĳi�S������=�m��I���d#�=u�h������!�����bC7���F�cƯa�(�=��w��}�n�W��*|��i,R8�� ���k4<�!Pv���5w��d5����cq��BT4��)u��-��X�eEC�p���\*���蓼!3P��k�^�H�ث~�P��2#�s�ZyO���js�xq��H�{V���x����u��8F�����c��H�?�)PNojF�W���5͍�D�x�~�E����/l|���x��X&2i��k�64�V;Z���q���`�ؕ
�i��-�X��B�li�bF�r�r	SM�G�0O�s�Vf���׹�-V Ż��yWj�%��a[�RƈL�k�XM~�ә�XF��_�Ki;�NGax]�n�l)�!7<SD	�d���}�E��QK�a7���ŵ
.+���>�oH��_w����&� �h� '�}���������qP���
��ѯ�����[�d`��Ud�WH���=g����W^w#Qu(8��Ք&��h��Q�枕<��������~���@��>�S?����Z�����;�+ÀF���]���toe04�����[�a&)L�̈́"����
5�-֠G�+f`+yf������q{��:���wڒ� �s|V�<|b���Rq�Ff�l�/
�7D����f	��i]�K�f�$�1Di��u}��A6��l�j���K�nM�i�QWչ]�}�{�v�����>�nd��O*��o��4�s��x��->=�f���-J
��/�L"�]�!���^�+��)=�?�8�Zl�˄	m2��:w$�A���C���:Ύ��o����J�(�p� �簜5H� 'H��X��K����C����}�3� ��\�_���3�t5��V�<	�&"�bL��6�n��y��z�Re#'k��� ����_�m��TR�F=6�7v�9���g��Ļj��%d�Qy)�
D^�_Ŏ������&�1���|y��5]�����(��e*��y�N�Z�$W�b�r	
�p�֬��M�+NA��Si�9f�*/hrΓՎz�C�L1���q�.@�]hNTUF}H�ֶ#���u\���&Lg^�#}�e�2��G)�ฅ"�*!_����t!0k��<s���}��ޥ��[���~���e%��8�+�^��,2�f��RJ�}đ��r+�����'/tA���_�Q��,��k�Я��]�&4J�v���E!��_�]}��S��I�@Fl�J�@�<�Z��_�m�����/ҩ��H�ۘ벑ț��;� ?��I��-^��'��'��
��a��nQ5�Le$ʿ�qE���&��e��̭nXs�8��P"p�.
��K�L�W#�03���:=%�BѲ�t?I��,����\`x�:�cv��@�V�g'��E��j Av��%d�������(�K"����*�tEOoq��U�?���_���� ��*�J�#�nߺg�ލH{�Y=�ە�̯�x�`�� �l�K jT�Z}�$|sn�;	?�΅�=�v*;D�3�?����kW\l`�S�3�^�*)���N��4Ͱ.��[/��q��>��{��[��A̛��@�AAzܞI��v%x�a�fx����c�2d��zP1�2^�L���6q��0�����<�m=�SO.ŉ�!Ԛ�����e�`��5�Ȋ�����])6!p��/ӎI�b��.��;>2+�#�1�OY��A�+;�囫G�Uץ�n�s�| i��|3�]�������^��VӺ��ۣ{�dVG%�^7ʋ���:]�?5��o���+���%�;c�EG����{7c{^{��u3y�(�:�Jr�6��I����@�������3�5DVQS~����*Z� a����Ip�>Ɏ><��3����a6l�!�Ȝ�kF�$w��c$g�*!���q�^�_e��Z6d���%J.G3�S�]E���6��$��ٮ��^Fm�o�ڀ�7�Q��4��P�ï��M_��6ҵP��7Ty��u+�3ryFVw#��p�M����Z,�r��2*�UF��
F��'�Y>i�9��O����4�p�J=�T��͑'J�I0�.���%�p/���v������e+0����(���7�A�H�ƽn�fŎ<��0@������`���n�z^��&�]��Z.�����}�,�q��r���Ίz\��+�ǜ$&֪�Q5�f��X��M,]���Eގ3���������-�esA�F��t.����U��'�]���s�>���5K���3$��*c������o_�ێ9�����r�F&^P��zHrr�,aҷ7�
9;��B.X�<�*�D�Y�5£Rt���K�M��ނ�ڕ������n�1H���P�����@���ۛ��j.���H��G�rx"Sa���ǈ��Q��������3]A����vҏR��Ҭ�0�Q��2Ŕ����0��ϵ&��N��Q�
\(Y��돭Jj�3�������或�H"�X�z[\�7*�ʍ�x���P-�>�2ˇ0(�F�h_0����2��Z�Y�2���.��H<g�����V'\ы���(J�0v�'��
���:TJ{$�\;E88�('����9$��!Uy�O�2d����I�gR���h�!����e���t*��'�k҆[%!1e�R� 3]0��gt)9K2�-��t�d3��Z��"/�]�0�4c[Ѡ��%FN�ǰ����c�^^a�2{�0Y�'
"(��^�Tl�l�}$�,�8�"=�"��ٚ�D� 7j4��NI���|C�Y�a9�A�T&���V�"�){��L�#����a��mB����Q������.i,q�_�#�D��jL������i���,��R��k�9,R=B5�m`�t���%'D�	���Z(r����B��l� E�/��\2D���Bv�O��,��5DX>��X�ձ���ZOJ7�.�aE�g�Eт���$��X���vLgR�9��z�o^���YQLbJQ
9K�Yb���������9qB͑�#_?�j!Z;�k���#.�f8�1�|%��KN��D��
?'s�����%d�Gp����F�A�C�b~*��SZ�FA���
�i�$b�3��CF�z�&
4�;4G�`�	��U��{�ލ>oG�*"�7�U�wV*pO�]z��F$SOᦢ@so�t+��o�vvG��%�s:t��y��&�}�(Ey,
vV�8K�{�
��x��}ed�|V��4i��b��Ӿ�?��k�����y|�[@�%�����1��J�n���rv�8�MŦk����}��:j+L`7��KbwRG3G���$������v<�� ����h���c'Աv�4���à�z[m��ϩ
�V�]e���V��r��~-3}*�L�����srm���y������x���?90e�:Z���\qq�߲�v���&�NeZ��vZ�(�"�? ���nc���˽�A�쇦)A��L6V�W�Ѳ�5�t���}<mF}��Hv��o.d���ⶠ:�8Z��s�^"=�]�4m>:+�
�O�\��O�D0����=�9�	3�g��Cs�n����&�����'D���{��	����HJ1^���F��$�Bg.Z,@!�9��^�� ���k�/��k����T�ⶈ>���@��h�Hk�>�˺� y�:�t$aIa�g� �ꡔ���� ӭBu�=��N%n��]��y��`��{���)���E{�w���@Z�u���&ŷ��k���� ��Z*��C���VPkw|>ω@�O��=��a+�\H��4n�Zd�Y�m��]'�#�Zu���=�t�
�Ր��
��E7t�ż��vw�۹�t�Z��_,���/�H)Ϻ��Cd���5�<�����F�87�}�Ⱥ[dҵ�!����Z��0z�D�M�gye�l�<*��?2%{[D0r�%bF��!�b/��;�w��u�\�V}�8�_���'���&{�i��I��#�>>�.7p��{R�"��q2��{��޷`{Bs�+��,�Y����.�vӧ�=n�8�D� �4�t�i��h�}>������ds���0���G�`�Vq��~�#+�5��i�`|���
�#��cV��0]irZ�[��C����f����ǞmY�&<���p����q�{�1��ܮ֦�cǲ�o'�O��1��ƴ�L�^�uА�(�?�LS�_�P���8���_ǚ��B[��E$�h6�YX�{"�y�����c���'u�������ֲ4;Q�+���wST�x�[!���p����+�K�Հ�7��_I��f��Ħ��g
���k�o��-o�np����h�m�h3�:D�t灕݃3�nL��� ��a6	��C��{ȉ����W�Q��������y��}������R��
i,He6��\������q"thK^$/�t��GE�C	��s'#���\մ�����M\sdt�}�X�qT��H���m�1�{�5^nk�8��2���XvE��(�^�Bx���w:i{�xI:s��hE�h���&�%i~��z ��4��RfMNA'砺�^�{{�P龾}yN��~��_���o f��������8��!��b���1}�A�\��۵	�W��W�_��zil��Ʉ�D�ΦI�*�x��{��U��[ ,�m_-+��E�Xc�.E�F91y0�T��p7M��"�o6eZ�X�b�����������?wY�%$��Ϧy]E��-��
�������[8��e���<"�c�E��N�U�*d0y.$��-��5�!k	 �m��C��}�F]���)�r��.��xFME���ȧe�7>(��f�r�B/�E/`��ǯAgXo��|J�M��f=�OM���W ��ti�},Glw�D>�i��&���KJ�eē��>���j�%(4���I���"�<ϯ�w�m߿���tN��K�UY@!:���ƫ�-H��9�c*a$��Y	��.�� s��'�U�3�� ��*O�'�����v���o �d?f_'ċ�aO<[G�k~V��|�ìA��������!ƽ��Ξ5�b�����G��k߈Fʺ=a��ZR6("OL�M_1����RI�OM)E,�������E��▢����7 ��a�ߩI��e�EX�=���_��Z��Pm���6��7]�jU?��w�fC�3�hrw['��։�EO�#o��W����MY�a���)�2�Ha���7�JF�����"����}�.�6A��w�b'�u�}laՓ��๧� W�싒���cư�;9ڼ�_�>�P�܌�����׉L�C쭾�΂��>NyӂG�Gzh :O�ȸ��Rrv�P�$5�dm&�^x]��]���7�[M��?_�����A��w/�k��D�D˿"{t��D���Bj���y�5���������#��p�SNb}�0#/��b�ᎴD�,�y�c�?.����������I��CD���Z�ȒN��-+�E�k~]���^U��"�'���ձ/�Ș��p8w5|�����Z��� ��1q_^f�90B�m8�~�iɄz;�>k�mOb�PNء�O�R'�u�Ypo0P�vh_�W��Of&���	�jl]�yۏ8�,%Г\�H<Ɩ�S^�D���k�8��1�a��3�.Y��fG�{�K���(����=�<^�[b�rݓ��(1�;m0��I3<�zݻ��NF�`�O�S����7[��ݢ�A|�9"h\I~��&�o��r1Ĕ�H����t�b-��Cɮ�߱0�S��7��?��I�}l�<��y���f���Í��fj
́�z�8���ɉ�����KȔ�_&$�{�(�G��w]�7�}�Sz��u���܍��6%�E,�,w�5f�r�ԉ�x��)ѬW�ê��u
hLP!���$V�����e��\m�$���Q��AR �)L�;��> �V�(P�1T�G��K����Y��30��^���RX�v���|l�߻a�jpĂ�1�e�ϟp�g����s@H�lF���N�Q�"�!���.�xS�tV���� x���r��r���^f�5:����H�%a�-��U�o��sP��|'ll�M;��.{�	�8��iOz&}ÀvhS/��L��.\q��2��
����\:����WMg��,l��K	e�*�L*w53�i�|)�Hi�V|ۗ�]�Ѐq���gSd�e��n	y�P�<Y�#������3�iƝ�yگg֗� ����{�E�³�X2�F�=��@`�(\��$���դ�_bɉ7@pg#/�٧��oy���p9�ki���=8D%����Y1��qA�,��	�$��S{Y����sn��;�^EW��I`��62�|���l��+��Ks�����8�=�	�%}S�g����ς3N�6�jg��a�
4°�e�{D�2���lW�_�Sl_V+�6�_)waj�[;��"��1\���1�K��#�]vkC���~M7�(�&�9���g���p�fۇ�Φ�W��I2a �p_�J�s�Oh��iM@~�z�oE�H��9+ �..��d?���þ�n��.�JQ�n#�}�D+�`zc���z�*@<��[� ���nڝJ�L���*d]�F�hs�pB���XV��7����kYK)��O)��	�ݱ��)����x�޵���k|��&Ia�:?��`cc#C��W��Щ���W���H��Q�/�$益��x��]*��)�U�Pk`��W�~4v-�VG�!�R�A���'�����_zbjQ^�)�Օjx�X�� w�R�}D[�2mcϫ��r]k�����r�@Ui�Z6���Qq�4�C�Sbγj{5e�&;9}[[;�=�����2	�Ȝ�jA��.�F-%��G|j�A$ͧ��E5��$�:+�;��������8_C��_���QP�o^v'VBoU��ù��I|b�YM#cm��A�>lâC��>lBx�G��;�m������z77���B��~�o���xk�ڷ�Nlx*Յ�ҥ|�A�Pң���T�t�RSM[���Dm��+�<Qi֢3��FHb���+�X[��������V��\�@'�S�V<؄�B_!�u��Q��3�����2�w�#�#�-*q�����S>o��`�} �`�ɭ�R�Z��g�C�c��T��N�R�)i��M�O��C��pJ|� G��3�˞P;j�X�ea�%wypg�P
wy���&1��qN<*��++��~ڷ�a)KF�t+V��d�%��b&�Ҩ-c�AֆB�s��L���gxȇJw���B�����pP����rR�KF$���:�����܅|63T 
�͏?<�ɵ�����Z�j. Fg��.�� ����#Bj�Rw�J���� $�BS��Y�q�:@���ZTh���� o�
 {��EJs����u3U����n'�<GJ!d�j��vvW��&�Lգ�ލ=��)��(M��"���ŪɆs˨�l�X�<kDw���|��K/�Y�$4Z�<����_�U�F�M"`0��qrր�~�c(���t�
���'P;d�a;� ��}�6r�Ndl�+4K\=�PX��$��F�CoP��핢T��sz���H��-xS~q�s�:ՆX���ǔH�f�	�H:��43�DA��a��S A�nr@������*�y>����@1��F� [&b�N�	,�;�,�ȵ�����_����_��--��Q�a$���E�����ڧ�ղ|��&��vA�aG��d< L��?C�k����?�KD���,�I�|����~è�U\�G��u�<�+��i��/� ?�.t�� S���jp��;F٣/
l������?�A�����$��sM,��H�E�{4Aa[�=1S5�l�7E�h���P�/u��%�}�$U��g�T�Dqx�ީJ��Q7Kbq�
�D�:�衜��r������+a��?�x�>����y�e�*.�>A�����_�pN#�j(UK����f��7��AYo�Eww��ݕ��	��}�/~�p��P=�爴`�/�xO�`<���6 ț�Q�{$`����)�h2�?�2�5�� *��sDr�)��t��T�[�r��z)�ꙸ�{�D���I�(�������l+�@S��'�xO2�/9�O@s�ݡ�`��J����=��t��Tu{%E�����&��}����=�~lፅ^�}d7�	@Y�A�b���YU6�F�޵���3dR�("G�'�Q��^�NeV���$c�x"jpɺrp�w���ٕM<"����v�H�yr�-O��$������ֻm�i��g6I�>���?c��q"2�2�0V��`N(߳�ƶ7���� ��Q`�	�J#�\ue��':�l�f��T�ْ����~N��>uE�]�b�
d�>��#��VH�Jz�8���]�1$�����Z.���8M�:O���8�s���f	ˡC"o��,�r�@$V�G 9di��5�iW&/)����2��0�@�6X��yG@�!h�NP��o��Z��c��q�
��l�,|-)���i��)E?�����[ES�)#����aaR����%:L>y��Pz��a/�4����~�k���� ����u)RI��A	]�0�����)ayj��|��z�F�,���V!j:� dtJ��>
��J���+��4�ܐ�5 0�ȷ��(u�7+nqz����x�%�1����G� ���E��ƷQ�PV�Ly߿Aya'A���g�1�o��*�D����ޥ��e�׸���K`���I�Vx��=d�_T~���jd�uύz��en�֛\�z��=J+�e��p֭��a��Ŗn���B"��������qEf�l��
���k��|>�$\\i-����	;�����?��4|	5:�t�Ӥr��#�8DX�-2���gy��Ri	�2�A:�m���x�I����k }*�����)�W��[��v#�DpM[F�J�'��{̰���yVW3�gh7F��y`�o?ڳ��/a}�%����J_�������;\l@���a��,��@X�OrW�$�����ӯ���?xntN_�p�F����7��|�5/7tH?r�ѷ�A�
ga�ʆ6��G�l{�}P5Өf?of3��O��W@�@>Dm+�����RYq��Va�8[3~c���ro���"<��|�R;�=I]G����;���l��C���0Q��N�lO�Q��+]!�V�A�n��|�����8i���~������@1HY���9�b��M7�e���8G�?l��6��[Ʈ�<5��"@�`W^
W0䠶>-O������/X)���L�|v �(k&����݌��b"W���
6��>�90@KXc��2��b�R򴤝�҆����ľ�Dh�9�g>�l������L5��a���|��f�!��
�x]��RŅ�ȎD�*2[�D��s�"�,�Ѯ-l#mr^�O�j�i��!+Iɘ�~[���ߖ���Lm-WjZ��1���]�L	���w��u�?�Y����To��/����lŘ�dD�
Vb���>��*�KT��3��"lj~u	aϹ�6Ѿ�5F3�vu/Se3M{�I�7A��;�z���]=?�����;T2B�V�j���zC� p�e�UB"FYK�>�c'%Z�s�����_C�]iw�ۺQ<s���}Gyħ&jM��90�o�+�g�z�C��Y�S����y����'���ܦ{��_0a!MǙ[\{'�t�e���a���15�R}0��=�ݿ��{hE��lF[m�&`�+�ҶV�
��k+q���q�ѩq��z�3�8�T�Nq��d��#�@����k��쇮�� �����K�Nh��0O�vF�e�)Ft�[� �h�4�v����%0�!����ė$�D<6�iU�`��x��	/�G��?&�+�C��T��t���Lڧ��Ш�zLå��'x�4��T8?P!F"��u�0���[�0]�%<������1͵Љ��(�HM�\BY+��/X�Q~C Z��	��� x�m�85�S������7Ax43����r3�&�큉!|?�Pb��@-��PTeBb�
����	!��vF<��u1�n�e� �����=�G/��L.����SCr� �_�0����ˑx��̔�.�4�Jw@n���*�F��=�n����Iw�[��_�UU�KaH���7�n�05��;4���Ν�OI����V"�x�;�(h��}��O��!��",g	/�fW�n��)�h�5"�/��V���j���tTa2����$��F
6���a��#��aP�@�{�@���M����y������k/;|jT���!�9j��3)3{S��X��Q��tY/������JhB&�-�	�1j�v�ffJ�ڼ
�������[+����8�L�/-��L>D݃���0dK5
�q�����������xx�8�N����/n���h.E2�vtJ�{q��.���F�ħT�JJי�Z>�-E�B���4m�d���Д�U.x��p��iP�hܿ�������ŝ�ӤC��@�7�<�`Dk�NKrv��ѩʰ��5C�4�I��ݔ�c�θ�7I�<�F��O5%N֯�� �`�$|5n�[������{�M�&�bpR|$�7d�j��]�sw�=���߁�o�(���r["F�a��[�r���UwmǞ�O-�O���c�v��$dK����;�U{��>�����n�o4P�����4�j�o�/����nx�N��h�#`hk�y��M��Ju;���� �+�˟��@��FS�x��V���G'hUۃ�L7Ԗ�k�7�q��&}*���O���?�ylZ�Oa4�h[3��*��ۙ=����������%kh9� ��Z�D٥�fJ�{C<��ʴ.�,�k!��j��ROF���}�K���8����wm��A�ej�Ɵ��`$Cu������ǉ��{τ�ک�ä1��H�����hL"�a�h�TD+��{�Y���9������f:�(.X䪜G���^2����\��Ԕ엃����HJ�Ne1� ܓ�^fco*Ȍf�t>vw6���0�V��9	��Z�\t�� �7�v��zbY�C�k�RUl�-�MB�n�e/�]��I�k �j��ySXYO�/�+c3�p��ۣ�Y>��Yc�-v�[jI�V&v#k�'`�o���|��r4
�B�)d��#o�D���ۤc `��:�	o)���B&���6V���/��OIO��Q���ӣ�a���4���'�q����z��u/�n?j˚���m����T��Gƪ�`fw���6Al<�#��@�'��J�%*����J����?n���f=5)�,�!MI�8%��ϋ;7������a7�j�M���^<9�`��<&+"��XB!g��a�(G�adI9�ؠ	-#b��	�6ͼJ{jg��Sd�N�Jl�L�����N)C��u��gE{q�Q2�q������-76��9�4vr����ڪ+[v�B�(9QR��Ed�aq��By�ܽN%os�pV�����l�x<�g刍��Y|����,SK9+�C��=}t�Ww;��\&I|ʞ�0��>WC>�㡓��|�w��
��e�S���IԙB�͑~�z1�n�a����k���ݟo1�]��RU�:�}
��Q����tBȥ'd]������K}$._Y��X	��.J��%�Ouyx��!"��*!
��ʉA[2y��
?�Q���H�"���!߄&d�2�D6.n�b2`��\����
/�����g�a�C���~>_K�������Y��GV�u&�a�Ih�Ȣ����Z%��~b�J�/�أ� [�K�\#l�M�W]��3ַ����xwY���u���e�v���*��})1�Q6�49rݧJΟH�G%!�G� �c8g�ּ˂�>b�&���������J2�������
"|�1�!���X?#	�����!`4̑4��6�./r��~$��jS��Edw��`��=N�n�S��O����C#���Q3�-`pZ�ĠCz�oA��x�p{m
.nGx�E`����|l&HE�)IH���ћX��9(b��,%LY��g�}�@�2����]Q�eίĺ	��%��Ը�Ѧ��Kwxd���(�8�BԂ���I�sKIS��NK&,��t��C16���*���aI�Qy]
���V+�`�rQ��ˎ�f��|�Ĝ���aa�����������c2[y�>l�b��zF��ܞ�v}�=A�|;��
x�[�[g�$��q?֣��}V���d�5c�?��-���a�#����z�� ���7�$��Ol�Z��/	P�n�a=�������aw��C{�5�Q/�np�;���>�9#�b�a(��Ǆ��X�{p��5`Ҭ��j��� �UY��ˉ�:'�\�� �@�K_!u��FF^Nߋ�n���b���0v��d�\�{�sEC��	ۄ�ݢG�/���_̧��EnVǲ�9\�f?TH�&�f���s*�,PW����=�E�O� ���7qQ���� �߷�O1�O��C�$�R\?��{�U�<�ݦy��
׈�U�ېF�����;�k3��q`Z�'�5�Lz�#��PY���X�	kd��p���Z�[���0V�������w�fwoPQT(<�y[���zk �J&Z{c�u�:��ƻ���(0Z���f�4C9��P�f7�ŷ�Y�PF�P{���_�2 M�����<�q�A��RWz1�]i��_ �<)i�	�h�� ݣD����s~�<�K�a�C�!��,e1~�ھ�
�?�ӠP�y`��q�՝��amP1e��]���4�`���� FD�6�o�W�v�O���>��<@�R�f[�n)P�߰2�IPC·�DW�a���%��F���q��CB� &Q{��-iM�f*U�+=Û���0f�/���V��w�c�K֚L'y�HR�05n��=▅㭂G?�7��FM�x-\2;�S�L@HG�:�5��[>m�f1�QL�y4J�h��T2Nԩ�5Zj���,{Z��֟Ah��8y��3<
�����j�k�x�4�����3��`����������Sm�%��b�mNa��
r�[��v��dT���@z��l8���@H���h,/>J*�i�s�:ݏ��tx�8����c 8����k�<a����.�T d�_.�')�h1=�>�g���bs�d�8�b,�q��[W �}���G�t#�c��q~���YS��|G;^���[��Gw8~�/c+�֑����a�d�r�������e�?f�B�;�B��������*��|��d��~Y�*��qu��N�`:��!RS�9Q{� q;�0f�����?OJ��)/��;��eE�U �E@N�dQl�/�\�<�k�c���;Ɯ>���wY>w=��%�K��`OSI��kW�ԧ��X���P��{�����`�Z��ø!�eD���`Z����rm��Ʃ��陶�U`O3S֘����̅t�f�����^��_[_�)�v}�F�&ǅS�WFjmh��xQ�u���R�-倐�v8R�hS���:��$�ί㭝&�J�C�Gŗ�Hd�#R���m���a_1!Z�E�L8���hf���@�����]�p��XW�Z#�79��;h�l�����f%�?̓C�yu��kͥ���%96΄W���\W�� ��F������ ��B9WLd�=jv!sV������YoE��G�n
�!^r~I�}�}���������K w�	��>r"}W���	��C��2k��tsIHo1�U���Sǣ'�����M��2�ڮՋÙ�ӌ8[c���旣.��p��ʒ�Q2�8�(�h��fC�!���n�	�!�Af���&�3Gt]�Ζ܇IO����.�
�lz�:�W�^�d�aٞ���q���E�Hپ׳��N��]j`��;o�m�h
#|7�m|B�خ�j�^����\{
�����oy�O�:�µ\��f�.^]}})����l��v���4r��Aց� �Z�r[M'f����t�+������8�
1B����5	Ջt�^%a�)�>�R�wɬ�C�;Xc���]��qȊc��
�j<G(����ʬp�Bҷ������㾋.��X�P"��n�Rc'�U���r0CT�?�Q�p0��d0D!���?��X9���b<�ht�
n���}/v��%�&r
���⿃�;�j\$we��<q4Ӹ��
�TEqYug�lj�7��a+�R}�����%ŗG�Y�72������,�B�W*�P���v��f�^�ޕ�g��f�	������z6Pfg��e�si�8g�u߾d���6�ӧ/-
�c�sK�.��'�b8�!嬏�2(a=���t-/%5��� +�Gz!L��s�H[����xB��˃��N��ʊB&��	1i�;��w��O��>qo#T��M+2D�$���t�T�س�Lݶs��9�3|�	��S^���0�?4f�}.=�߱�fO�F~w��Z��� ��`�VX��3y�%�����M�t�d�f���C�i��o�5����#*\z+B�C9�!l~��Z�k�ΔP/�g9
�%q]�,�����^f�Tps�dv�vw6׊�:4��ѭ���ƅ����q>Y՗�+��B\���p��"�����e�/�΍Z�vWx�.� ��|�n?����dn�x&h��;qy�Z�����zC���RoY3���b��p֭&J���j�+�
8#�Ѫ��$��E�	m�%C@W�#?�b���]]@3�[����4��X?��Ҕ�/�׼�2�lh�P_��.��<���I����+�>(�A"&���~����<}X�I+=楜!1Tc�Ov��5�U�]:I�a�K���E	_;���7]����^���m<�!K���D�Oq;�g��/&���tq��k�ls�lX����!�i�8j�'�=q�[1ꭼ�;�hvA|VW���k��N���M�O���9�hػ�7��U���l���.<�+5�+�/���#�꽼�~S,W���@�|j�9�]��*8����QI�*���
�W B�`�G�m^�h:�%'�*#��[j�]��ֱ���i�Wm��ߝJ��/|Y�*X�vp5��o��^s4����ғO(d�`J/7�4 �D;��A��E�-�k��ӟ`?>2ɝp`2��2���X	���4\^2�O��6x�My�>��䃴D+�CU��oPِ��ԣ��Z{��7R��K��f��x�D''>�{xb\��2���&�m�N�ct߳��<7)��cȀ uc�SDאi�MR:Vq8#2n�,d3P}�}OiYf�Xs�u6b��M\���MP<rY��Ks~�)2�����DDN]����"�.���BKPM�e;�1�bp.eP[�?�$��_�;Pf�]n� �ec�d��� ~:tT��0��9]ޘ=�s&�-j>B{mX5S2{��~S��������J_���*��y{C�7��(���ϱ�5���}��u@4���+���dG?N7�ѫC^E�F�
�QOc9/�4�/�o������4=4k�8h�+���fl�m�A��<�1�4��ہ7�<���#␇<�bXN�Yʅ�EDcu{��wS��WM�E�_�'�������Aݜ�Xm�tӟ����:2H��v>�O�-�ث���Ls�e�A�e�W�\ �\w����,H������
���i����<��I����\l��DC"to�²�����5��\q�S�g��r�!�.�ё�l�֕�캆��TQrv4�o+�t<�ܞ?� Շ�RYw�cv����<<&��H���%��Om�׻�n�C��uO���OzT�S�ÆZ�%.@j.�����cZ��x��|ٰ7^RV�UW(y���O��R�7��Z�Hإ� �W������k������t�k���X䨄ڌ<����y��@�G�J5��%��O/�4�G�G�m�=Ψ�t���xp������:;�1�Cc �}��ٔ ��I=�9a�s6~&>4�����ow�ڪ۟�t=21���Ot�L�d��.�� �6{r���n|*'9�!�!1�TA+J+�_������6"Ӻ���X���Ej%l
�~��	i�6lc�I��q���_ZI�b+$U¸*B6'/�а���E�o���$df�a��Yo�#��#oة56[����v!�1����xĒ��Û��:��g,���π��1�J�Fp4s7W(�^G2Jb��Fs�����[���40[a� ����A!� @���Ե����f�-A�/�"�M��2>�ê�0��{|Q�ǵ�R�����x �7��c�+�#\�"{�,{�l�r����s�c�0v�XlA��9u��篿�j:�
1�-��	N���Ccl��W�V_�T>Xyt�Ӝ�~
�/�~`�N�*�n���o�+��'���0�
^��G,�"Toc�����݉���RK׈5�u\/����tq@[�)cr�����~M����v'�
B��iRM�1�A��e����f�w���U;���}�0�$�����r)!yF_����������I�d���[���8>7�H}�i.4S��tfs2�
�)i��/��y;��a����~{*7=�j_%��Ĕ lXDQn���ۓ���6��#�gZ��1����e��kqb�3��Ѣ�����|��Lj�o�7r�ZB��6P2'�<\�������%�o�o�Z
�2�2�i#2�%}-NBd�*RR���'X�
b���̾
�.�Qg	������	�8�4��ѥV�h~s�%�ϩBL�5�o����)HK��i�e����0.T�U#VB��M)���i@��}��񵱇A�H�>M�P����~�I�z@����c��M5!^��}$��b��.a[���80�?M�c-������qquJr�O���C1KW���2H'#c������Zh�:��j�Rs��H�2��5�ߜH?�#�����LD�}�{U�J�ZZ�� |�D2��#Tr���v0����c�-/L���E����i�)�A�<�DZf�nRKKF�ޮcT��+`���.�A�ȉ���b@�7{�QUr�ׯ
*�"`�������	�v����4-xՍ^�4���$�%A��5,1J��b��5*\�)� �����{��bWt�g�I���d�O���ڀ@³�{*���$�������QօU�;�<�	3�汼���U��bB]ј&}p����Li\�|��0q��m��ERlD�c��Z���G|硗ψ}a��9�;�-�/�%�e�/;#�4H���QbQ�Jz�}�r�����e��>��g�%@(�{e���y�3��qɡ�F�A�]H��9{=/��I:�҂_��o4}@�ɾ��?�[����7� Rk�T����l���Jiw���d%X 0��e0?��v1�V+������hd��" 6��y�D�|M�3d�s��6y�7�-�eJZ�w�p5���ݣ��)o)�� ��z�6|�P|MB�x�%�Buܿ��U|\��*xd�h����`�:Y�VK*C;�{>h�6k�+[�>�_�Zp\eS�^��´J)�)�t��̮�ZU����l��aXg4���-� ��-PZ��>�vj��ZX[����FUޜC�"	̰5���ʯdW����-�-��ȫЯ������53�sPФ�9׳*��7�3���K3
H;��@Ͽ=�>Wg�Ut�k����A�/��[&n�����Լ���h�Sh�54T����vXV[�T�/�|zP��cۇ�A�6� ���5 N�>���S��h�d���9�~G�,�-������ ����Fj�cY���<i��Z9�����X�'����s�T��ڛy���O�Չ�HSi?ɂTֈ�������	M��y���0x�KvA�}ݛ
�lqX�CF\�q���kPL�~�8����X��R�֨V}��G0e����!߉<UTc5��tH:�LT~���hd$���
4b륆��7K4�D��~^�p��:���O�`{Ҫ�mU؜Y+;�Gz%j|~�Fa�p{��:�qB\jM~�OK;����ы�v�w,�5��WD��Ӎu�"D�pb���������K梴K�K�n��b������d�l��s�\�P�Rn����tbp����,�ɵ�.��$������f��J��h�� ����k4��4�p��I��3��y��IZ��}w՜ L7�e��OP{���m�$˳]X�j�l�Pd���C�7�����!�n1w����{�
�<Q]ԆdF��5;�9�bVR;���W<� "z���[7c�/2�0E�o܅���S�U��t�S}`��H���V�̕���e�b�r�W)�p ��w\�ɅÁJn��/'Y�eƼGt4�2�*���45k+�]�;����I62�`}�/��Q�1��8閶���g�x#3v�% ���VO���O�k..N�r�������L���gJ#��d1C��"�뽻X�8������0rV6�^43�I-ˑ�!J��M�'ɦ�����q�.'��Sh��8�����v3�Y��
�8 �]+IC1QW̳���Q�ҏ�r�������]]t����`H�P�!�(���+�~Q(Ӿ-RՎ�t�Xuk��h��/�`hU�[,$[Q�/����T�XeHȠZ��8���+�Ә�~#G���I��Э�X`�Z����/Z�ٵ����S��@���x=�b婈Jr���R��a���-��AZ�{�.7l�[mq@�{G|�Yk'b��}�l`C�,j&��g����q@��N�o�|g���I�˒O���CX/^:2F6x���s 7���ȠJ�a@b��ݰ�i�)Zr�b�p�ȟ�V�o���9qו�]�̰��1�5�'�,�0���a,>'��0|#5�Ǚ[
�
H�Ą��h����_�% �7a1���~��`&�i�.s�9��o���&�.��33jP��������f.]�7�hE���rH(co>Go�MA�=��[��g��K�B���68W�P4����5Vӯ|�x�$o	?��<�R�;�-����/���O��opg.5[�x8�0�ﾗ�R�o�����+"l���a��'�t�y�{����M��j�Z���-->A2���ll����#HK������~B��<Y��	7Z��i14��K�x\���圆ZW2C��8��g�����1�տ�CE�./<�K+�Z�A�ܛm��#��/XV:Ǆu�zF_Cѷ���PǷM��*9�vQ�k�ӟ���W�,^d��Wހ�U�-�8Jy�׸	�)�-��@ �i���e�<i����ii���ݶ=N��u<ݮe���p��9ү�h�j����(�1��� �ۧ�	��qə���|wq��H�u�Zk�Q-������՘ڕl���R5��P3�5���/���k�$n�y�R���7Xf���:�W�f�7v*7�����,���X������bHr�v7ɽ���Գٙf��:]��!�����9jv��4R���"U=���맡�X��I鬠Y�o�F?J�U�FGZZ9�`Dk=k���dM�
��K.G��ęs>8�bW#���d=�.u3DA��`,��� 2)-lύC���>P/�4�d��5�_�,��#L4`^�<�R���Ɗ��ڊ�6"��iu�j	��7S�a��o�Vs�����d�=�T4�^�}�_��Kea&��x�2E�6:^��d*�:��Q1�K`��'����}�|{�jp��������wd:w��K釦�p5;`N�.�_f������e^����_?���,l���e��7�R�=�W�)�þ��?�0�O���2gS7E	bA���#���Ǝ�ײ6G����v�פ�J�-{���p�u{�@t�"��q����U '���Y�~F,jm�� {��$�k ��>Ѡ��D����*�?(�i��_0n4>s�Ȑ��9&q�G\a��xBƌq�@@3l%q,�>�L�����G��c�_W7IT&��'g"C� Juo���1�0 ^��i����>���A�5;~���*K�7;0�З&�����l��wׄ�^Oi�/��;�rX`R���sI�����ɜ�����%{4ߍj�z�!���Mx]S��Ƣ�~>��$�?]E�ع����,��2qR��?A�Y$U���@�JD�f��|Gmc��N𮎰����-1���3�㤎��:���L]AFWp�t��1�I� ]����p�gp��U�B�29"���_%��la0{;��<F���ԑ���\�ǘ���}}]Y�p����Q���,z��k���J�6��d�a��D6-������C�1��+��b;�9�`5�L[G~���T�{5�褢�K"4��Y���|�D֗�>�Y�#��T���M<�)qCp%�T$���\d:7;��0�篽��+U����#�22�� 5qtU�X���=z+;�����xcF��0 �o+E+s�~�!<�װ�W��TL��Qи�!�w��R��UEр��	���!�&ʜ��"g�F��"����+g�5 �������w1pMs�T��Iݦb�WQ�ݮ�b�t�m��yM�����z'IVz9t�2�_�EAR���=��.HL�/�X����
�1����"ԝ"��L�aaϸi�RA��|4Ǭ�'c�d�PcB|��@�d�M�*�Ѝm^��CD?�_&��+M�3ؑ�\�N�L
��ȟ�!.bI׋˹��X��5ɰ����_�<�Pd[��(=еsA�E����n E���[E]�G�&1���*d�6x��->�I�B��F><=��cf�k��C�6Ԫ�k¸�q<�Vc������򖵜m/�>K1�P݆�#���qA��3g�8\�`	��n  �e�-���(+��&S�\��l�N��Ųd���g[�,�	��o�A`L
���>W���#��3�I��:��0���p�����ź��.�`� Bڃt��i���k����v��>��cNރF��%��n���"�e�X0�9���w棱��<3�����o1'5{I<qs$�Y�p��X��(�d�Ac����V�쭫E���|�1v��Z��D�Qy �j�0�7��;jk���!.!!�.[dV�Ia�P<�W�M��m��b���$�_"�y'9,��K�r��+�:&�[�P�er����
��ĩ4wg� �������+��NCN�M_�~x���+-U�����vc�YrZ�/�\ຎˡ�Vu��+��$'\aI�,!�8��V���D8o4�pD��F����A�w��n�bY~����2e���M�x��U92ő��i1W�ś�,��LJ*�M(�(/om�x�_
�DV��?����s�=8�ޝzǽTҿ�e[#"&{����5�mj
���!�C�Fp�U�s܁n��k����7�rIA)KB�����y��\.���o1��e�C��K��уŮ�^�[�[>�d��{0�֜������� ��xJ8>��� �=����E8���^u�V\��C)���,��j�\�N0#��Ij[�t�����Z}ʣP��ESL�(��a���E\�lB?D�mV�D�%���ǓF�/U�9����8ͬ���"���n�0��P�G(��Q1�(t2-8Q��A�ɲQpڈ`$zX��d5�x}Ds{N�q��_P��T�Lk�m��7ޱ�~��1\9�p`E���2m�-��n�A�Bu�*J�2��?ǘF��?;˩~q1ѻbe(L��כǼ �?�d�k����E�R���U0W��u%=L�NN���Ȇ�L�9�ӷ }���==d�����8�Ⱥ��;J�B�:&��L�����I�em��%�ۘd79G�0[8� �{���(�1����N�����9��O�&ה��ǐe�A�ܖ��©L}�����V��UD��[a@���撬_�� w��O"��_�xCز�$ V�k/�*��S$�c�����ℷ8���[�H(ag
�q���sK�:�H�t�uz~�㚤lĀ�M(0գa��|�U|D��TF����Rh�?X�Cf�sk�K��W�Ū�
��Q�nx/J�g}E�5&M�ih�Ŝ�.���A�޳w���Y����~��l�^�&?t4U�Ss�����͜�\q[莃Q�9�ҕڜ�\ H��J�|+�����&?]��wp��M���}��{.���E~�;�o��,oBܚ`tԐ�h�s.ba�ʁ3�7��ΩP��?~��
0/��y�f��%��Lݴ�:V�AZ�<=��[?te''�T��b!�[�.��9�o�و+rt��˳ �v�榫)�,4�|���� ����sV���.�Ks��ʸGk؏�*��S����:>�8���<e��v�gb]/�=m��ֿ����B�V1�PFs
�[���]����*$Q��!����|�U-eĠ�^#|�ҝP.Xy=7� )���k�U�}u�Ri��v~ A>v��e
���Dex�Њ�v��I[ +������I�Ţ��2]_i�t�!�B����n���uR\���6D۟��9�ª�H�R�dd�������5�e�S!GA�h$��P�����04܇���j�5}��j/V�<KR�eĢ�Cܟ�oj�H��C[_8bu%L��[^7NH�}�:���v<3\�k]K�L�[�/k�~�ީ��G��a���R�U=���)u�h�D���ѧ��&��
ɹH�[4�מk��w)*& /�MN�,����S�X2\CAEu��9x\^�h6*J���>A�,-��1p������D�ů���t-�2[��(�(7p��7�P�\�.�I hɄU��pm[��+��$�p��A.;�mf�t���B�ť^��m!��e���.��S%�~A.g�H�&���xY�6�`s".A�#'4��ua�����ou�^�A�ښݜG���/���ыf3�I>���W	�,��]�8,�������9�5�����5�`ș��a��1z��j	۰E�<֔�a�=N,�d��z����S�8���Tь��'a��K�V��(�S�}�[�q(����^���Д�Ҳxr���E�t�u�~�$�Q�Y�M�~�/�u�Y*�1���*7�9�3�ڇ��Ľ9�nf��0�W0F��x_��X�B_���j��Y��I�<.R[�~��7���>��}P���*�]��:�����Ƣv"�B(�2?`(��C�UBQ>���e�`�����|�LY���grD܆'-��9-��#�Or܁����_�Ѣ(��K�P)��!�_]w-�\TD�bI�U�Ɂq�s$��Tu3�e_���C���<�'@W�;��V��|@��� ��T�3�MZ!���`.�_��#]�F ������ٹ�	5T�����Y
�b�	��!f�u���"ac ���qɛk�u+���_ث+,�o��M,���k�;?sq�������o�Ld�_Z=�f7;��U�z��W���`��"�{�dڋ�L�	PN�q@�����+�~�y `mjj���D���{C�XzGT���D��	Q|���(�q0w�N�]tu�o���h��:�E��C�o��PrX�kd@	Z�L�x	��ԕ��ך����_�W-p��%<G��9�9�*��-�I*�Z���2c��!�f��R����-��x���p���D2�Vdu�n��mVvr'���v sgN1f	!qV���]��?W�>Vn�����j�D�L!S�S�	 �[�����1�$0���#\�� ;/%"��,��r������d58�f�I��=�|�^�GB��ͳ���?D_J�JJj�U��[2��R ��kQ�59������n�ڙ�3e��O���9�{��I���"��yK���P�fu�����Fê摤|�8U��Q���B��B�a�GRae_O%�!M�k�z�<&ݶ2����M�ȗ�-w�"�/<��'}w���\�h�f���v�p�/i1;�#n�?ӟ���b��2����*!��FG��S�#�!F�/��۟��ԫ(9t�>��]NWɀ�\����h���?���(�2e���=E'4Y�]7��w~E�
�j�����j87R�P�Z���Ns�~0��a�|6ٰH�@/�.�o��r���4@�|���m�G=WW��W7S�.v?�4�H�Z^r��(�[�����2�v�;��ؑ �d&NX�<���k�g�ҹБ1��x�̡d����fD;��PT�=w2��P��+��頽���(��v0;�x�>t�^��J<�h��й�E�+�^DN[Z2�\���%O.��R���� ���l�SI��XBC���������e�ؙ�i�דtD~Qj��1����.9JJͺ�:SZ3l%��+������=;I����<��[�jj��=�~(U*��q�4���*�TU螓W����2��L[g�51�I����A��H��k���|�KP:��Q�B$~K੎�,�DeVc�X��D���tꞝ-Qz�Df���<ɈLJ bD�:,�!R�:�]A%B_D��a�B����(R,�G�����̟p���R0 n�|��t����Ѡ����53�m���\6�p=B��4u%|�P�`.�����Beڡc�߽�ڌ�Ei�E�de2�b��IҀY|�x��u��a)F$��ra�.�ݢ�^M�t��H��X�vJ�_u/-P�����2:G_�y�)8�[�"j�PP��4̼"< `�:"���]�?����5��Ѽ�;{�XA��o�[d�w�le�Xi�!�qNG������F�rCO�1�4(|�+����0e��hp=�fB����.xc�W�]��߂�|?dpyӦ��_��J��U��X��h:�C1a��T����K��N�s����h%��g��'Z��ܶB]؞ s�\���Ӎ�x&+���|��nv(�3�*	�g����	��_�3�<)�`j�1����^��L/�J���
��T[E��t�i嚕�����NmΉb.΀Ϩ��8��|�JP�迎֗g8zLݨ7,Ӳ@��TP� � �H}�%��>�p��|���0��'�3
?Nr��]&9����-���00�������C�����"k��)��"ӵ��91��S�>�z1K��8�ҕ��{EQۇ+������@���2���u�k��غ �w�:�����GP�F,r��uce1vz_󲥕 ��������	7W�����Q]#fu�d2��5��v��Mv40�hJ���Z�3U�+��;K�C�٭��j[�Z���JV|C+�%�&DR�I�:�V�I?Զ/����G��/�^&8D�54�@�:�����rC��D��/�d��I�T�_�0}3����?k��O_������n���eD�N��%);����O`�ɬ��g�E���N�Jj���8��A�3��)zaKރ��l��.��99�Sv���ɮ�%�����������H�A�F��}编�C�8p�
avJ�[5�/�{1����`!2���;n�5t�/s��}�~��Kd�h�*-��,��(��[���*0pn�a��R�XN���c����'Z��8����/��cX�upk�"�i�Eic�>�)"]E2r�)�:RqY>��oG)�'���)�� _
G���M2�"�q�!�!�NxP���O���W����K�Ɇpc�a3T���UA��3V
���n�#Y�*s׸\�B�f"�b�0���Ui����~R�-�Hm@�6�h���z����v������^�5�_�� � *�ZA"=J�˂�h���>r�ޡ�J�V(.ԙ�5'\��ȹu�N�
�{M��h��g���/�#?���N}�F���ro���q�?r�ӫ?i���ET @���NJ��~�n-��uR��MQ�ǟ���R� & ����ڤj4�O�vh�����]4Xgh�'93qv�i%e�R��j�]-kS��Y���q��a�ay���6%�`Uȸ"�f��\�X{����ᕩ�V5��#�4gi�:]X8��yE�5�Ӿ,�r�����$F9�u"�Ɉ֌~� ��)j#������@V��K�\�I��P�(���y�ţ�9����&���*��(j��S��1]흓��FR�ujy�{)�����|aꋾ�N�Mn�f:_����r�"�3�ns���_�Am��G�ʃ���6'=�Уc9���5�e��<�=�IC�ڀZ�Mcs4�8 ��5�D�jdC�%Y(���1{l�Q��Ԣd͔����";y�ɻ�
��Z�g�3M@�u/�m�8�y]X-B?/��2*}���.p�\0��F;	u��a������+�(�5����0�t~yK�Dn�<�a'�Џ,���+��f��l�p����w�F�d��S��D��(�;��.�b�dk���X?�E��f���S���k������a����!��X��a(�#�LS��TjI4�밹��U�-�sG�I�w��י�!ذ���1�J�N���Q�#��w�7CI�̚�C�_��gEF����~r-X�9s�'N�kI*�Ty���0n��w�].67@�ަ��Y;H>i�7�8~�����q�4m�[��Ū�&ѱ+����U�ї �l�h�y�k���N$,$3[0�Ss�	�Y3�\�k�mZ�,�V(C@��`�f�GXAdL�B��� ,`\Z0����N������*q;^�^��x�__����� ��3��B�=(軒��Bu��pg�r�sp\r�����{!g��?Ҫ��;\�~�Z����3��"��3����v��?�}<�٠�H��ĴF/&�������ԑ@X�]�<"��G'�GN�i�}4M����9:��3�&a؞\y��Cۋ��%ɲf��x�����A�[lAPF���$�^��g<,�����F��hN��q7�Yot��+�<w���䏓SRA�DČ0�X�1�o��0*����*ӂha�rx3iSM���I�x�-���~�kkО 8�:�+�wP8��H��Ѹn�_B�h�b�׍S�ʵHS�x�_��{ �s�q䋞����{��K	6���*�`Ə���r�0���ep���o��.z!Ԓ�Y�;
��}.A�F�#��'���xCv�������5�zi^�:=ۨ`ã�X�@��㍯ׁ����S��V�L~&�B@Ȯ*_3Wc�uP��8��C���8�;q�mW�����*k�I��a��mv#4�����<�(k��)�n'�=_?�8�h��N�ϙ�)�>z�;=�K�)V��Љ"��50�	9J�$1A����_��(d�5(8J�m���OY�s�Z}���]�/n�ݝ���aD%ym��mf����'��o�U7flm���@��_�i�H�Rza`=gz&��&�,� v"r����7��N�ђ���9�q��� �;�ς�'�c��.{7/V�z�g�W��(���֐G�M�l�~E���[����0|8�f�ߤn�uW	�ث������ʖ������tK;�jdg*�@Z�eF�'�f�	�2�)C1X�O��cV )���m�x2Hl�D��D��z���Pz�k;�5�:֯Z��L��ыM�i�~qڗ�tG�*,�%?��c��$0�6n�\���3US��U���}��i�X?ϵ����=
�g����ӊns��/Q"�@)�0��8��Z��;�^Z�����E7z,$J�8�X��������N�$fL�b6͆������wxGΣWFu��V�{�Xf�tP��1	�e%�n2��Ns��i�Lk�V�����|�B�o�X-�1�̆?�gm�IFѪ/f�Orc�H���u�rj&#,���
��r��d�����W����bFP&��eL���'�K�S� AS�����4hf6bС�JT?U�U�~���T������@ &��̄��rзCԻh$���<klp���o���xyS�]P6�S>��M���+��i����/?�b�S�r�B�9ț�'4�F+XJ5\���uqw�)qع��;�#8Y֚�EAD֨�KD��� 0u"INk���_��#�F�G�N�)�)��*��\���7M�V~^#�c������`�����e�����獒�˦�v���o1��bUԜ���.����y�e2�r�W�Z�Z�ݔ�%U;b0�eVZ���Z3{Q��;3�����x#��JX�v�/���Y0�:��T�#�v��QS�\F��E����9�XfZ6��5b�g���0}5�K%�Z��^�U���l�3�7��Y��-�F�@^�2*��y)�/���$e��P�"�lj��a��;kbŊ�q����0��<*�B��E'Z6��&�IG��w/�����%Q�qٸuY
i�x+x1�f����4{I1����D�)��z�lq���ׁJ�]Pس��9
���U��iU���*j��9�`1�k���"��|��2�++p�v��z���z�e����a�!��e���:�~�����q���o�2c�q����a�Ħ��].���e���~$�2�S�Y\�H<�`k�*�)] ԭ�ص�|ֺ��o2A�6�k����Pg_����g#��ܣ�`�	�E���ҳ���P_��J��^K9�b\��_�`�Ц�������ȕ�l�US��Ղ?�i}8i:&��5���Ю�L鯓��\Q�Z)Q�	I,B��dwjT)х���V�\)8��#� ��|�/���o�-~)�1�e�$Q�I/ຜd�;��2�N�A�,��qx�y�}�Wϩ�,Ve㿃��c��d�ȓД���ҜʜLkj��~�%_>Bd���y\�����u�0ׅ�8������`  ެt���4hA�Yش�]-{�~ξ��	͖4�}�)�5TDP�#��КT;AB�o�3�]��UU[?�6΢�q�������uK��2
;8�B�򄰼q�+�3���u�<}�Ņ`U�ץqʬ�d8���km�,d˂���wҙBc��"��G'm0]]��J�{��S�1=M���5ҭ*��w���-Л�1�/�{��r�����[��6&�4�i<�7���549;r�~��g��͑�'��r&�B�Q�k8�h�O7������[ӷ����X/�{���2'-�#ҏ���|�͈�)��pP�'~i~8:"k�|�^��B/�U�Y�Q�1I����3�{wڃ�*�;�)#uL�oi�Sқ=+�	�U���O����Xh^�pd��&Q�����v�D1� ��b���O���B�J7׫��S_�1YQ|~�N�}�nmF�]�J�g�sǏ�T(��\\H)\�unT���\��l�^"d�)��t��d㈑;oCܨ����V�G0�/͹!�2d ���\�� �k�4[_	�'+�t�z߯ �P�ǔ�>s3�Q�r�Q.=�/���J�`m׫�CY����V�x
j���a�$q�6;M#�`�"�KmS
%����ɞ�j����a>�b��v꿦��λ�ׄ��yڭ}����=fI����0��U[S�4�S���6�׍Ž����?� �4}߶�O�]6:I��	�:1 ����&�^�x���ͨ%�g�>�Lk���w��?5��5��*"��=��
��-G������>�&��ԓ��H����G,��+a�o�t_��F����q��w�#�:(�L�X����
_�5������vN�F�6j�עsF�n�q(`��s�t����ƃg��z���@�1���!���>�jB�H�hs�8��<�$~��ǥ�P�>*��,'hBG�V��}�y����{&"��-b���D��}�$��u�#���ꈸ
��u�������ahI=��-J\���K8
"��Ġ���f,+���r�?o6��f��-���-�|��
GIG_����y{�)����,��q������YU�p1y<�'j�k���U]�}�C��ĥ��&آc�mA_5!��'���̈́U�؋0���s�Y;��R���V>���upb������5:�g�4E �\�*b>Zq6?�Z�_p`�֜�?䞵��hO�{Ҭ�a��y��U�(�L1��)�$A.�U���D�eR��>s�w�=jSv����xu�$L����<,��k�u��?�O���$)i�j�fe�΁7��^��_�]ܬ8�ԧ��Ԁ�6>�}eq.�tϴHo)=�}�Z���(��?�~�3d��W)���;��<rA���Fe�{@iQ��y��e�u�ⴜ�c޻4�621���4p6L#F��'��Y���ɞ�=�]B�jJ�\k�����,����Q��X��觰���?c�9t�/?�Q�����l�^�b�?�I���ѥ.�6�*�u�BN�7���ѯ�< q��4�I���^S���������w�K��;"�<[��Umn��BY����AM���� >���BYH%ع�g�Cd�T�����M��5�hw���Ͻ�^t����������b|6zB�p*�5J�V�g�;ZMźbCY*+kX���"�]%ʱ�m3k�حY0#I�6�$�ܑyG����_���~}��Wq��Me�?�r~Y�Q���BN���t�is����\�3t�z̓�%o���	��c6�GcVH`�����Ơ��{�$4]�#��1��*��Ͷ�v�b@FI������[��w��u�j�)�۞r�")��ش�*����[J���yS�м+f�"+��&��f�jڔ/r�\�H��G$_\{^Go5�hP���,%iU ��"�c�Z�X]����ȋ䂩�[N��1ږG噀̍)�����i�猸Ӳ#��l}��S~4� o�X~�G1i:�~C�}V�~8�l��6K�6��T6�Κ�3��d�_����[u����.�_Q�#ޡ�1�33�����H<��3�H�*�