-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Bay4yXjDNbl+i6DlNxWPAVQdlHDBg4IpBIEZolBdER1C1+HA7gseGTTJ+lhF7esOaSl6g2PLdZmX
GK7/tU/AJzZDtu/yjO6cOeJlZaxgSD8etGsW4ZTphYR33Cr1PbS+Gwbkipv1WBm3fVyb/I0cOcAD
8V+E8idIs3NqeUSxHci2LO3o5gigNM8euI1JGgzoV9rubgtkDNTIXDyGY6+bTAXqjAkHdh/0v+Nm
xDc5JZy7e18od7pQlb+V6dEYqh8fl4VHn3OcXePhwHAfwjlib2oM2l6yvjB2AErptxGN3l9b5+HO
hVlksV0OXajOHgaCgS8LiwdKBpCH1MhNUhJK3Q==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 32928)
`protect data_block
SG10MgbVb6ytCfKDbczGF2Tw3OrdU9gzhgUgxAQG85izlU2qiwzRVX+r+tVT6Gqdg3+0wZe2ykRd
GPgy3F97aakfMk7o9KuOwZ994Eq/KMeF/DNjJ/H1K6QfsqW5mmKC8/VJ8JcnsyBme298ZFDRw43x
SJs/wl56UkbWk3mV9smhLLB+eiAZkBHu2J2b8lHBaieLV0nMccouSyi6x3Le720Z2rtUl/unQEuf
3kFoFzsoJ9VA0Mr4Ke5SQt/iKrB8Wa+NwGZlhwrfhPrUUES9YPWOoCoEpHge+GXNfLmIVICr3Az6
EE0Bj0wsMJO1PB0+9QZyEXhL+mTsHSWg1JcWnlcgEUy8RVE2JcOlrhYHstw+NSO4TIQWkFa+17WS
QyGm80MR9/uVvKDFPoBdOIMRvBb+3Q4Zl+g+uPZ8fx8cwYxTL/tFwE5LFFJaBUuPWM/VUS3wbq1f
lD5XCS8faPaI6gTzFdLNDg2fgDx+Tm6EMBzs1r7cygJ6cqyS2tBMGkVkXYmkKPVR800jvo1hWsIJ
RP8z9X3cAfi9+xI3k4oMbaJupTy/j4r++kfG0HL1/zlIFaHU4V2U/liGaP8RssuAyWCr/vjGSqNw
N1ynP8Rcld7Emznd7p0EzLkeEWwYdvbB+rF5tjKWUY3o84Tkjnz/gCxnZj35lsenWHy4sy/YRRxZ
GtG6MHfv2Ae6MFrYjOCm/tM246nfL5nQ3/TS7Q6kZKl+WFxAQ0MZDg+FHkQ2A3YCJFOhqyjKjUio
+wifGSRTC/TfDbyQOEz0WHbQPD5ZNQrH+wARIC3EGaKVKGHXtKqVuCW8nV4mmrBjd5D5ws1ujyLO
hUFRf/Ap60CUgmG75mPhm7zmaNERqyUeZckM4jkwRo4MHD3gBVcfNdYh458+lOsUddVeLA1GWWpw
j7Ug7EkPX5useHDCxnOUz4pbcetjpSYLtxP0OyfCYXYnTp7MccS1CKpooNyNxQtxumBnZTeGj1cw
ZcBqb4DoPYOlcnKCcd35kI1tGpNRSuRKOKpkZ8D18h2sWZTaBbHCtDa0p5q4f2DO3AaR9hUrvOAK
ysxkHywMM8wxs+E0UBwZ3o+pGuwnt90ssFxYunqgWBTZ1SNRdfzl4quApP37Q3VSCkD1oZQ8+fYz
fGPHnbjDzukh79A4rMwckHZgFq/wwv3ET4Cf4EVlx9PRdfCU9N1r7f6TWcGx7ZUDXEjLhs7mmG8V
uPdB59VIGBmdahv3Dl2J126Lqh712EpziiAB3CCEakqGoXg+VpvmULO13YUoElADKGfTEuTyzSgN
Z5onXjvfXol/1RsxbalTV4402xmML9abxiylmMNmtJ5H8nyqxsfuKkuNxA69CDiFAfm6vPu9dORk
rWZyU2dImHJJ5Bt0zMQO0B9gv93sdYSaX5EYvNj9HZVv5jtwzLuIrg3cICKluFCuAQC3DnyP/93V
FOlfAAZ0P/FNp83vJmVqr2ejgzZ7vD9PsVZ4AfObGARYl5HJlt+cKwbfvjuoA9x1QPLShOjnAMdW
I3AP7mmRy4avXw57YbMoB6hw8fg/IYsrU5Ckxk3v8EuDvsmwB6bfXq9g/DMXSDtV2RNhV4CFK0/O
dLsjDOUsGUPEDExibU+Jjpikz3Wu2LY9vgWsqMFwY+EIYtnooGwEFmvmm2U7GgEwfQI7xhM3MFL1
kHVQBIeTJepIs2SGnn1/492ru2Djrzd6YqxDKRG3Tf/7CPdMoAXyiVlT/tot0AnYLQio1EsL5Q60
F6DW+tsx7h0VEmYCJ6ERG55XF5Wo7tIL6ktYLRpgDY3HScb1gssfWiT0UG8NOhiG9WwksOPe0dBl
lXOCpPWgVqxgxj56Diru8K9bf3J/Aa9jpg6HEjstRGDLHvxbctRrFAGIeo6OsBFT08PMOQ6JbX7R
A+OeG7wygpLJBptr45/YDljzNRCtD4XGMRCUtJvhgn1nQGvZoN1fICl4wnGmYX5F3n7ySSB12j6M
3Vsoi3ex4pEz9qmhxZ1QhoyoQM7FbS5k3LRkt/2/wr4dZmNl9mKp5Sft4ZivKLdjGH3zTasWPi7k
teyRKdVqybvUmED1/VoyHedMQS6nIv8EoDthAffoQAs/cT+W2phx1778ws11flDs5/YxPykIcTbI
Srrnn5cvPFgP8KjImGJ3knoown/dMVHJ+240NR6WstszCs19RTG01vk7LEpieTkuEGtL4a+XqUfs
fQW2fJWO3ekzNZzvW3yGPWP7A0MoJIIl/l9gHCIsVuiqoOo+TyJb3U2dYiP62YzIYGsD2VNBz3bE
F3wRo5gOyCfeMpM2BPO2RwONr03Tv8tiNK47/uHb4f4h+DON/jv8T4h0qsRzmA29ZTph+0HrDXjn
XLdFlJsH57Okdn6zKO2geSXFeLEr7DLUhIGjUCXjMuQu47n6W/T1bC7kMwIKpE9RGzx5VGZVjcGQ
axOF5lZ3SNNXULJqftUWhrLY8IqsbX++EAhUSAoeGS2daMwK6xfE3nFVdHEIHFJt5IC63iZ5/Ug5
hQ2p1Wnd2AvAe2jHev/ddWwKaNnj2VH6dPNwi1j6fbQZl6KJNtwIkzvyNHHAbiKjE8Cll3mvy9+9
Zr6brds8sSkktcyZOpw6rp6dHSVvJ3lzEcs4TQZrVP/p69TbucGEBiomkGA/v+0dB8ZgfVV0JEYB
/tcLfXxYfSrwKTwPyjxCiQp/qv+zPS7PDZVHRXK7wNrELu03NbgCfCltQ7VTfxB5cCmE2KmprF31
Pf/p6EywB0i8as6DC8E+EakpvteGhbWe5AWBeGZmHezmIm1D6PrA79S6ljX+EhoWxghBuBM6SvJK
XhnIfsdg8WQoqJ+JSHKbZl7zhjHqQwogsJPyW8m62p1CX+1avIqqU649KZJBQ4YbCUMAZJVPdWZ6
B9/VsVamquEt96o6TygkSI7NB3FNvDDEreWN9umGGo9yyQ5fMH8ZsBvPYPU68roFaZKJujJPX+pP
YUkk12UcMLkG9aU6eeQ4Ync++XuAfEFaQTAaxAiOCFleMH73jtxP7K45e8jMpiQBiPUJ2I5AUZDa
91tlOUuDbGUC224DRKjsk6m8pTMyTCFuEndSxd/6+2kHCLzh9bueIm6Gadq/WgZaJLeQ6g7JFDm0
kE3GOmXlGjv0AIqn1DytuGDlg0PyHSCU/BEGc87dfh+Ojoblxun5qTO0rzLZ+ALukURUopD6WOgJ
UDyJ28P9oAXB73Noe5Gp0yVf+6YoNGLLzSOf7h/e0VY7vahoX+2FY6ZiWwTBXV4eGYrt1FVsNSX0
KZhuss2FId4OTonhCYvQHAQ4RS73tWRAQbxSw300LTloIGb/IMY/Oxt5mGwVcdl0lWnfiwxoxGuA
8CGhIUx3chz6IBLgX0ieTAZt2jyoyHHRF7BFZ3KpqZkX2I+3JD4+E4jRT6FHVnt9syPfj809z8hP
V6Hf6CWOkELZIY52SpqeRKwJbr2uHfJMLqyBNjXyykamLtEA0WChCsmFmdh4cjTZjfQVe+HizLbZ
pzTHqKcMTNOsAAPzNPogWyVv7rPE9dE5AesIz3nDXlJVwAvyWsAlvJiCgEfd+IRk8pIMXsstk/5O
cPbBhiKpBDzNAoEy2qibVTFwyx2OHJUc7Zg5dVSZBttPZuOn/zK3PiGX0dFkLXO0lEy+kZOC0paZ
162fo3JiJRTGnHxpqR+mX8e0Mm9bf6+j7LNEJpr05KivOjZ3fdZ5l+BE9vgN4JQxM12rZofhAmLr
QuJ7Thl2RylOAGu3z4csIfsfSlIoDOhCu0158eQV4jRpCpvM0+jm+8uViEqSKTnNTlJ5g4vIq49g
aRa4RPvfCGsXfOzCgPODHHxKyzhWSy2/DtEpyocxBUjo3s6q7mOOzPOZi1E9rZBdQJ4iIL0YP/W/
M1pgRho7ciaP5uFoIhTuiSsDKDWWjPBNf70PWsjkWSzjOUZO+N7fs7Abuminf0IESiR/YIcNE209
e64F5+UKHtfcULEyJWOT4zhyIU017Des2n7awQzBX5I/LB6DY6OhJ9uD48TAPnN3jC3+RriWZ5o7
xiPkwa0LjIBcD3JkR/47e/tTbr1UM76qbM2a1rFFs4LFRSsOSNCTfUUUcKJNmCE4eJ79LT4x1m+2
QOy0ObGNRxTEQRYcBelguIrowXqfRZxiUa7IMXUeNdrZ5csPFZJ6tEIdwtBuWY7nMNnImx4d6LJ9
vB/cD0r+zqLgSkyFZ4vJZKBNxC3fG1gigSGRrPvQIgC6VOIcN3bb5BAqh53E8HGa0mv3pouf9Wzn
DrFsxxxbcESYJ8VYarSj8S6jeiYDfM3eo6n1SiZb6/8BZro9wdZpnpxaNVQvjhQNxa03JmJ9h5PD
hk7TLZJs9lQ1SFBTRYBdUEd7FCiN+sOSdaob4edN6yOt1kqMCMrWi/5M39V6xeDjVVSurx6pE1A1
F/5c/iaJekeR4qbd2QJLwPWZ2GYVgT4ZREPOvVi9DxekFCgN1J40LXUBsQUcXi5OpAWP9Mo14wF3
CoGoYdnzbktYAs0GWF8lVIBC8wQ+iwRAlf5pCTtEOjKAl2lrNOZkfSMYg4cb9qDUc8O3m1b1tYvq
j6QQrgyXNXu6nRcDJFiVagJE33liw0G3HJShgy8E5GDXsisYgytW7MPqRnCjwrPnYYuElJ9iFbbK
mba8QserqocyVxk1W8uPEAw8yPYILxkrnAjs/+HZBaXdotKr9ST3DTF//Rarbz2tkn6gYjv1jrPr
/gZNBdEzb2BBNqR+ZF8h2aPg77CctT2mUc+K3oaUzpGDM42TNGTB7e9/CzEZmSaD40eFiOZ9imUc
ctaYRq8NsgapdzHOqMNbahZJUkyC52uSzUy3FI45cTTxY99kZ/L+CJHCK8JRd/sCXiOJ1F3T0qZE
fbjesRqOKDcQ/C0AnMN/2kiB4Xfv5KOqngZv6nP9ZlXmmvUl7uRUok4NDikTVpnXfDQ6ZwHFiwSP
SOQ8aFCluwNp8WhNQy2AGMBRKfl+uoQQulhlRjWTydx9QxJmnM13qp1RPCL+a5fNnX1S3hb84fdh
UGJ7pElGJcvAZjZPsqKat27hoqHZXeFO3ST+IuIUKjI7f4XDcqjxcjS1BqzMrOMhN6qJSBAiuUD9
iToDBezVRTtCDWRzAlKSoEoEoxX1oQTWbHDLG3HJg6YUresugcgkEnlSKpSr52GpJIxiP4JNFu9k
QYHwvtJUUDZiWHzwRChy97DbPlV3BX9GJcZeMwPPmj4Vra7tY7MBxAkZY5K7UbPkrMd2shKLYAZv
hmIgxQXID2+DUnNETY34L3DvMPmEkk2k1CSn+G2HC0iufco2GSJLWQUEyp+KYBy9DI+rzrJNfiIh
oY8f4N/OF0XM6rfHVX83vaLjNWavzitCcgvokO3ULJ9/PQdxxVNTf15Qa8plbIOgM+uCmXYBT+Fk
qYZlsFSz1yLLmp3g+CuD7MUyQjADpj6R6sRDDDSgD2RN79+Aq66OfSxhKr4HAE9J/5sK03O6gA8B
MGQR6Vggf/wwSXwFT6Yv54y6CZBIgWn9By+ny6VfZNUBVjoMTVOcwChSXjsFexeeu1xMuIyGE8cf
4av0MHPIIyhrWraID3NyD0kxrueVSm6oi3s+AItAGcjaOkqn8ULmnTH8yinJtfZ+6AlG2NoE/vaJ
hF415q1f0qCQ0Pwg9RYNM7V4zo801VMuQVZ2oQVvkY/44Kqs6De/WRordGFo33l3u25ZYs14bH40
dGK8uVuUfSvTfpHtABAQS5NcVVkJp5RhrAw7H5Iy9Id2c22X6ysrdcIS8E4RPnmGEEHeDovZHFy9
dsYifYTB/EQHDb2/Bh+1XlIYj2sFzp3PLHFGF6eXmoe+ItxMj+ChK+/mzhFsrlayLVPFBQHNptbh
jgs+d6UpAbOZCXbozEBvvnYPNcZRzopRTcxdOUc0BDQyypYFMqxXGEU5nDEuSBumdqMmAE9NfMfS
sb/+PR6nvqMspHwFNAYJNuUhYebnn0Pkj5EjR5mLPrutxwgONyfwr+NvcPuwFVEkYMRKMRQKG9d0
Xv2yWCnDCR4u6D6m3Q1+Oab3M+Z9l2NsWnlicb6UNB1GkKJb0t+mYeFXpxDGAXECncDTrGp4YVlD
NGLzH328NdTbJuo20l5LbtmuAnjN1sBrY5AfbyYhDDATlGkllmfmTlpxFyyc1FUl9pxhqI5gsGEk
ATtsX70cezXcXgyHi33pDc9V0LWKldTDNETAf/zIyX/WVOINHs2w2aak+Dch4QZawB3fCPMdHxjT
Q/hmIjPZzr3FBiizw4nYPZQAQo0hJ5k7vtb03LLP28jpLmEw6FaulUstsGV1d7MyDNgDbC+KWsaF
IqS7PbLTsJ0xZrDyr1OysSKdxWmc/Ve7amZPW3RQHlEG2xRgzRxpHQdRYUktcqts0wV0/qW61EpE
UfwvcpYrcdAE19sIukG4Y0++lpDk3uvRtey7eRittG3+2KT9JhgBR1Uu2zOJMsZ33xpiFc7L6MRy
MRezhVeMzNjgrgk5nUxDNK5RQKHDZFuHhZIw2Y2VGOgLAtN9xobBuDz+K83Fm3yw1iDE7s37XIY4
G/LFzdEsqSIf4SP1IVEytc8jrLEwBtuts3qPq95kKo4RHQcIEF/E/tnLLe6kGn5g6tOXgHWHvG7T
pmEEVfpP/A/vBVGl8IMHVDuRDukvbLLM8YVwakSceE0eqEsyaPc9zn3R+l3ADcBhFvqmztARRx1O
k3ouDCnP+j9pXQp89QGT2VPuMxx/tZRczqu4D4t3JFOMTvBMNTFF7q2osKa6qAbN0XUt0JUYnwN5
d2HZD6ICLjm5EX0y9QI8fUNEL5LynzCD2+lPycD6QO7POC+0WRP6Q36QzZKudWNLTnm+jq3J86Ur
fDlMpeXvB+beHIF1w/OfQhYhcjDiMDttN/BOeS0PRuTrwHVx9lTRELyhtrewn8Vt46fKf1hWKLG0
cPTCwa08XOe/+mFw4w7qFKCXGlrvMcOAho+TFaC7gQtNO9fsu0OfmZzbk9BY+JiQhFcYsVQlbMyi
QLyEj0pUxhPT/XeUeWxCXzwVLB6gCrbzJvgCzQLoocA/OTgt+2LFv/x6pga8juLOnP64NyVFOnnp
gTrkIScBSDPfJPR4jjQFMlquhquqlyz8EkMaRJlPet7zoh3iQFRTEmTHdFhjzX2Ml//4d/kmIx7U
s25B0CLDREqvSmSVDbVB/SMYg3rW7Ot+34tQb4pcLf0k4i9RC2kUj/gxlqvvbZMk478jFuK/YWpm
T4ZoThZ9OvWqSvkqIkP8qVwl6GWbh8iIywEEphbaMz6U4ZlMnJb44WnClvkcboNtQEGr+3bd+59o
wtI6uXJlAYPyHaXE5H22TlaY1i0cMFCbvEplV55GI2oT2NGdBqRBjX2rVIYvJtYRbGeg9AAL2BoW
+R3N7MJtuJ1THYiORVDFPBGu0Afc0OgGeHDenAI1IsxUJv3qqzUcuEep9WF1uq+SN2cYZXdIC1oM
tzr/JlYdikq0ZybQmex8LJEhld/brZdBMYuPcUvKC1WJBmwhqIQHsYnWWTtlky8zT9dY1t9OryVC
VtGJQp55NxXMpPab3xcw1KLf9uz6fNESJaup/m6ZbLEzV0Pg5falap8NQVmYwiMF7yI7hW2DU6y0
+u+SEqOWQLo5MqHfopXrgnVJr1lczXUDpf30QP4z+JRCa7lddq5vLJYGCgdIqtmckWVjZU+Fgjpb
dFF0WIuKYpVP7WQC4fs2TQncDCjBuKlKhDV20kc9WcgAx8fF8vHVV1Xu52IFTIv8mJqgz4WNCKkt
A2Q7eN5yuRxiu2Ez7xWZcnoFXFMTNBQv4TmZWV9zTEfvPx4QF6VBBKq62sMbJ06EqjwWy2sn28CW
/Bc9oIzrqCLXmWHUDdy87CKUxn8L8rHBzJS9gKKQZnl7ePyvWoRit7SKpRyuc45uu8Q4r3F9zJ3K
rHJIvKY46tYq4ZYTxRfAD5w3q2X8cpGJ4A+4RToMhiDGs2CJK1fkFBFYfF4kn1R+iaUnv+J0QjqL
Dne/UVjn+NrqP2Q6rCGGF30Q9dhiWGFQ0zRAcGjOQ7/S9Y4/aKI237fbNflv5sb0hUHhXuBWr4Zk
jn9/vY2Mxo5MbvETAT/xArf4EHUnazGDGY6jwmaQpB9ELf+hfAgtLvF5baoodMtbx4b3k6scBmc2
pvQMQb+UQmvsHCKkDSbJB60ywhwr35rm9sbvpaOGNBB+OcZuId4REJGGQD8f8Rb8+8buqqlIiBgf
6Wld/981W6WwxGqCYd6o4zXDifv72fVbQbC5Okg9BqJCbZ6FVS+43ld1i1FQJdtW0bUqBkVd3QPG
jkxVaY2DEVpD0DLIor3QlQoAfGdRp6Ec4QbLPgZ8TSuX5kppFYsRGx0jAi+7fKrNgQhnth5C6DFm
fzmNHelXuRGKHvIrjxJAv7npwgbBTb0xelK1jN0I3xej1aFRrh5KA3vgtDhICKGugSv/0Dl/xG4S
hli69SIl7qorojmXhz2AfDrwhpTJcnI/t76jO9t2RLSI5HNr3cJa+yjq1vz8elYfeuq/rxCGW0v9
Dl8NUeEEbfPTAcOkc6RopoYCzJ/A6HglejUMG1AU1xw7ylONGP0ZeoVDimspu7oepdd6nMEanjMz
cJLS5zynRgk/UFCb6osaRPGtXHD4at0L/RicrBljVsnvrnRybi+zuOnXTBm3fDh0JddNcMwl+58i
gCFsCbBMrvKD6FXbsP/EsVP1icfsMUOex/SvaNGgo1WG4cq+AyqW/CZQ6W4lMF6gbHuAx7ShBCNl
hzG4Td9tHU0Ct/v1AOUaFD6T5/LAGoy6naKP8TGJSMQ/xwNiyO+JDCcFVvg7qDfJVT5q6vz1YHnv
xxSzfHRrfaI7viRs/D+unR2oAkmBFd1k5GgKsfEKtYP8I7+Fmi1YZ7zkU61I+suC92o+t7VTm/tm
x7BkpSlPSGe0xwACTmDzLviw8cq/7FwBnW4oX95TNvl5yk1z7W5tQJWCCw4uCNrjquX51Bibwr3R
wsEnOcQ2MKFV/yvgNt/boT290KQiKFxs/AZa3pn0q1Ob8FVYmg7hYyYLE084THCxqMGTX4XJzSPZ
TAFR4bju3bUTM6Bvj0W056F0V5AlRfbtTovkR8MWwx8dJdEXK+soW6r4F8E/kxZbb/LDhPjt7ZA9
znNd+/8GfzodUydW8gzhYtAvI4yAuEbZfjYWLFnqeDEPC8ebCn4g+BamdJO9Dwj0q8R8E8px47Gt
XKRB5yjHT0f1ovoELostXB38lSQl+nNZfHN1mmp1ocSnAyTw4uyXn6SJ8V+lrJy7kSpAcRauVoI1
nSq2x3heDvqY8GOGwsP2+TNSmMjqXgiXr3won6211epvm0HUUa2I5N1jppPSkVfwt9f+ufG4b95m
7ns+wJIA+1Aacr0nFryFJsjfPsNBi+Gut56M2GZBstni49T0+Rfhk2zkveGHINKX/xp3iQ2n3XXC
CAgIpkAx1CGsf78NZ8RKfA05MSOOnEwNvM9YvzPHqnFQsQKiadMl+4emZqGTiU/5nSam3YbUhyVn
RbKVBGBZJ16blo46NrOktzdYa65IFfaH32HCJ5Wk50WTmhsUJ1W0mOLXMgFvjNmetqKaH4mWJftN
eE1Nn1XdZKjATIIcIL74O+IsJBGxrDXvclYgNtvNXSCoErbe5ecHmgRPcIhaiMmSIEQyk+gd4lS9
iGtFDt/NItx6tiPIvixWApNaGwY/C8SjszJI2eZhe/0uuWMe4bxa7OgcaYF5T2tv4n4iKMXN0dGT
gfXD3H3vBKIqrSiXEYKNJBHIZOO9ekZJvpm6IYUb4RfOmFx3QNs2flyWDD6qF8dDN8/4EbN5vKWr
84/zfx4YwskoE3Sl4LBHTQPWtIVy6XBYGpAKNi6H/YGIi9M387nBxgb2DgV3T2rRU186AKzGIXES
+/HcJk2Bq4Xwenh59uCQuwms5fxsmLCuk2FhdQZnA6w4bfn9dedWUo87h1hhc8F7JooqjdcL70vJ
1OhgucrRg0zoXtKlMHOd/5ZYJGY28EeiZzb+UItoREK3lbMylch2kv6b8uK/7ucYDbYyW6hxFwRc
ZPhVgxm7425pkbzJWAuYH3djBimJw9oiNQuE3UyOudjtdd9f4mYFHRqBOxH/TZPsnmAgPBpkLPHO
KtaEuFzwn0niFPBieebQ2Q4BETx6gmJtx/Dv/Z0hSMiUUcd2MV/KFhkEs2Ws8P7cIEhU6y5kuwUW
1whYrGQnaJOYwn2CoO1ocUSushf2gkBUdP4pYbRSmvv7/Qjnix9gs4bvkEa3t2OBbaNoRfk/+a1e
1NUi7IrcEPR2Yy9zbTmzZ7eL6dD6mgCWYEb9L25Gf4pmxGWIjFIKo3RIPEUfWphP774Vz8HK+Xs0
CTLYaAeMQ8fsSGkYpM01pwrvhbK7mBE0VTUWaqRvlF9Fs/ln6k1r+v5BDSTQyrdWTMop6KzyA91h
/Q74mbqBfu8xaemI9vXqKTLj17LkDR4OHWvpCxj3CCMZ9VZM70ceSPNENJZBmuIMG9hai4ScGuiy
kyIgeqBybFzeVFkBWqw4bUXf/+yb+lCYX094fFfXCv8qidubfn5bvp9+LCs0WHY8iS7znpP3uMYi
uE8x9piClnufFI62zuJkk5VXEb8d/JycV+00T8jpJ/kGCnj3C6TyKg1FCbv78o5ZWdseWIyU7Vnc
Im5souKhW24dScaXWC2T2R7e6d5F0OhS51O8ezNRQMJeWzbyKWRYCaQnzEjQNnVumWclH9TNxMly
SiGsXo3i2skAPBsN9FtlHtpMeXWl1Oj/4XhlBCGg8Wlf0B39sb4dafbFY469F60kSQnsMHo0ll8i
ec9Ihgb05VvX3hCPQfQy4Cc2/xGr7RSi4+Idc8FPilvlwaDjb5dscPcPVH5b6OyPKoQX2s20/I+t
5m2RZrhzbqhNXtWgzmS8rQByt9iGelZ4yEOeub3IimZ8gJsyTQt5D0rdN5t4jPTV7tuOL6SLXrQm
C+Z3NHt2M46HSSMX5AffgiOkityd8JtfOC6nQ6ZTT5wIzuv6ErWN18gOQboW0pmyfM9IOMIWUNUx
tQ+wp1pnDbF7Wyk4xhJu8r+pvadBe4PejF79wXa1oyC3p37LkiuP5NsAfXFJ4zs/uM6hftTMU9Hq
Q7VEvnnXVsO/wopflgydPVd970GCW33Ryzz/p5uuwmfPW3txeM+3YtE5HCEAUgQsCXwQKjZxcKpL
oBG+qqo/dtLdwqmEoaDcg9QME+hSrVVJJrqF2Z//feiqp3JKl1IsV3PO2oLrTv5k0rAoiPXkVIas
ncQcXYOOyXeQgUnLagxfxxYRIEVJvv4hDNuBO4T/tfQPLQnmXOlkpmo/IrxnymrG9QP9TfnjfeYY
sQ+wumnwy2TUAUxgWhOOpO9Q5ZwWWSVlQxxmrPcjqk/5csolL4hpqvM8pvuz0N1kSQQLA2O0sXZn
vb2eSbiAAECg03ibgk1S+cUb/vGHmJ/Gp6I/woPk5FRE2Qd27XLJEs43SC3o/eOTglMec7pqPQ/h
OgSUcgqAvetq1M3Tk9F4L96Ijp5+Rfhqw+9J6EqiukvCUInGMu4CvDmX0o2tBg/hsnyeiaykaLo1
BCm015IywZ0YoJ8eHZrrWaCLVQwMbPYMLJHLsVzhxJxtGdJs7T2ip8WbHV6ZjkUzWuzFK+pdu/q5
73xoDJdwbUpxXjLAtLu2mE4s0tjtXr831FfVD+U7keH8fc9wdSlw5XfuXKFtqZvrX21StMVcPPnk
eyHq46+P34tUGw6taOJCxggZZbY32309PXPBmnPj3pZV8Aht2Rc8got44A0LCSVrH/4oJPmp3b1y
6ChXZIueX1UETRf58V0mrIu0Zn6/BSNByFK+Fv7LYd7xqysZwyyKVUQqnyEpTBEEnT1Bz9Qfs+ri
ypRznaaKsy6ulppa7dGFysghB4aFHzj6p3x/ZO9lUlTWQUwzNy3E6LBn7Enp/q/WF9FhFLRQzPiq
q6C6hjnBp14RXyQQGShoEg9sM6D+v9iMceDxs0iZSFL/5w1D3mpgp0+PnBRogHm8M3sqSYZ0ubWr
IO5Td8yeO/Jbjg6XjUvUqxliIhpMAT+PvWXHJbS9B4A9NOql1uGoTEgH3pdK49mEOdnkWKLsN4r0
otSJ3A62QpVMzZgPdqFUYWVNwSd59cYHIFpbvCCwMAvzhhZElldfPE35CyWEwe9JdSXQIu6M1Ajg
Iz3mQyavKJk1J9+QC8g7He7KTy/X3Vqlq09g6HB01b0tXhCsqx/nKlRXpHDcOxOacZPPHsmdlTAl
qVCDlv45J5Bq4PGK1QFjuyZop92NvAk18qTQisVmbWbh3Y6RPkhy9t+LVVvuzJkYE1qRRaSBVFEt
4k8u+Taj4XJJHYP40AD1iJmhHV5tW5yH5fltKX79xNB8nGz38VUXJh1EcNbFTz/T7e8A2tqFrmS+
eA7r4ZVirc8jfxlRMq37KZfo4CNPIEZ3GoQoNfIh2w/6pisXc4DHgdAXKfUACqBcRMIbPdG4Xvva
+08LteX3XPFvOF7JT1cFD21SFn0m116q+LZSkNRRR6i/eCqxuNjuHDaLzm8tqryvvH9aNoyD8tSp
dm4PIWXJ7Tb7yh7vu5ZTOjkQbeBGs/LPhRde3Mvj/fZfifDJAS+DDmNORnAXUqZ/mT0mubEzUl9t
i6/35sqIvnxhFECHE3l1jX4Uqszc2yauGE/blDsVZOdLnqybzbGREaHbStQOcC8UoLNDatrjI8F3
bsHf9YGB7GUz0xveiMOcSzlp+9aMsejSGJyKB7md7SjoPdD5kUZQNNCiwO8M7pGDoeoy6vmx5hgQ
JfBOqerhuSUIagY+MQFuC9w/l0wSxizFhVUvTPF9fsbFWRNJaHrDVt8NphsgUs8UVL82tSqzLoC7
4fxSptDHBlLLnOW4+6NhT73SIcyiiKpwIwgsef5wdRocCaRP6CKe256q7t2r30JpSQCsIg1Jx1mQ
bo5mXaVb0QuEZVSRGFvLgA4VzVHUrvkUc+0LJvCylFTvZ9hw8idoLGxo6ag8VvUrX5hZSYpl58Wh
GDQ/2jMbaBd4AOqQhgChsu1hjocCKJfrZMoMny/dtazrZouTLJIcKSEp8phqBo/yCkqsqxJI7cSC
cbf9j4pZk3OB+6VAlwMFiQPpDOsdhHWC0Jp/IGvgGodO+YdAi9n9mw4dccyX3s86QoaxBOBda+vv
MF4nBDCvXxMGGMGosUtHLEAOxoD4jKPLU9Nkfiq8RinHY+M3K1gA4xI6lb0wYMNNtbdn7aujSDPv
IqwVqbMk+F+Xvb4JRF+g/SvnFeHYiXR1QQx+S+djTSWj9cqZG/h82yhDSD+ATe7CVlaybC7UOJpw
xbZ6wbzuXJ9WMMfcOXEtrib0kVNbXdZkyAoxEm/6A0d1oZrTvrHC59n/uLthld2RX4xOZyoIWvM6
q72TNLne+0MVvJt3oVLaC2qJgNjOwndNW0UlqllJrA2tF+eQfPc5yazyU8EEibcQSqlh2oNy5Jkz
y6cXc22Iatik7tXieC9dNNRXAMV2L7O4SHRS7u1kBs87J9ZQKenqx6bu+uZoCSoEnZYJjl6QG+lL
Y6wWkPRm/x7XXhlXfgRcGaPa889hTl2Qa3UBL0V+qkGDM7yYe/OptpL7U1Y2l2WHzcOU1qw+7YSD
dDI/nxlQCwu9q+aSBclFsTq9YG8tSHLToLFk9HmyXSLAaMoMnbml8tKR47Yot5Vg25Q9RGGVY+AC
xdECreKKnewlUnRY9Nu5r/f4f/RJiY5pQhIucs02rSaFipBevzbNXJMp9oZ1fL1gL8nnfW0FfTXj
5P+Xb+kalFPyNuyq8RRZsFvxB+2fRLj9y4CIwAk/AJtNLIHjmfo7+oDH5esYb9iE0Iw0WqWMYdMI
A92ZEzqyPyjkwb6exxgzBFtvijKSR85UUPdq0ZmnGnuV3YQg+ZSong4Hsq54U31mnNe5rEqdKrOI
zgcd0BbxvxRDR/Xep244aayyVUKUFEGFsqP9xv6iEXSGEJLgt1foWzSyn7TWG1/HVLi8+DZ5aFGG
0dFtLH4IkB3B/mHKE8ZDLBBdB8wCLJrMWH3FZwtChkSDpZZ/6FQ1C/NjZrdffoqC/1Sf0QOdZaGk
bJSlwAK7JjYOcU6rdQhXRHPq7AaR9EkG/hshlchB3CAearAz6b+gXo9f7+/8rY/wZ8J8rL91nsLr
s1OAkQwi22Oj9xZfB/5Bj9hZkO+UoUeosqWk9GFCOQMDPnUuGdV3IMv8D6f77N1Pr139aVjMs+j1
xHBMvfU1wvW/W8nPNIGOeqxfJ5yQqLfCJRYIh+pCLZfg+AfMV3aBrntkLwZUF+YtTthzBDbmB2dP
nF77riwgbIoL5qkA3f/1l1yJ9V/nRIpGyXUBQAHtCp2B0zvalw7cyRDyOi7Pk8tzdV72R1HjiCik
9lietn2I0pRW1XfVkhUyg1HGHjKyU9G4ti6GDQdTf0gsN/6N8mXxGciyI+Iqjqb3+M4AfOlIW16Q
koPYCN9wwB2sNDq2fsQD5nLGJAfzwexwNh/bPjpfBG93lCe7CZ+kM+PwSjFKIjqzw8/w4pIoCD6X
lUmfifesebGT+3ZNda7vXSUIf6V9wKUFbXEeTY2NqWm1g0aFvbE14RfWEWCJW/5Ayvqz/YcfPd4A
Kdgq+qsRORWSFHS4UvMHyWXCVtUjLnztgpiTHGQrrOoU5Y8Xp8PycvOwV2tlKEQbvSvQn7JM5HNB
XzKog0/IqNjIa2SSgtnDux7aySkL4lmi7kZ9sQQPcZCNCn8eif7rLC6fpsXmYP4GSa3/TTi7N0mD
XNXGxGJ1ObNUtOYSUgIb7VCeBmybPIepURZ86UT/EYHddn64f8JIjA1Q4ZWe6FxrkRJ0JSRWP4b3
9q97QUAMsuxGSPZydQfLGAfDjCo9DbYqe2dKlEPIvc66YyNn5V9CVLZL7zzTcxDuJZ9ZfRSQJFc2
5cAsHhqXIqIiaei0CEkESkGlnyhrwrqC3+Xu+1gYJ1C8gQUSS23wE0jw8T3np3LwBlAtmglQrk1+
dzQQzq+r8iZIvLaGzSSelm3LHnqAGwdmHUzmD0Kuk4mvJEM5oLOYrl2enx4OyLLOGLPkmzw19Jvi
7yqdEvWS4PEhB3gGwfwC9HGPELTMOOtxwfFHSfC5NFQYs97u3slqQd2nAcXCp9UPIaVXSUOfodlc
ICl9nWSpCjq89Ug+KJybO6QSAayr3uJnfXJCBS93sshq2QJJRDJRxGYMaX2QvobAD9zTapW54xM9
MYn0Mq34E4Km1FOYYlrRLzBwiEcdG+CD4W00UL3wI7/MfdFIEMOYD2JmTvl+GVi4PBipQYrV4UeJ
3zmv3m5KdlzGEy5RITviTg9+P/qWFCcwI37/JC9LZk8bvcK+rInn/R5hViabfEepeNIcWgdd49a7
oBAqkuPblyS2/bwCtGEBrDVnja1qtOQj3HBHMMhsxNI39T8fqFUHrqLAGffzeRk9vjAYlhdY/Owf
ktG+KGtuegKfIIiYOr1I+paZFzW2t86i12SDTwyykNxvzwPw/hQ5gZnmyuazPPZnxVv3k0EAtYi+
iRKBxODtH1+ralV3isWtq9kjXHhb4/A4JdyNearTV94mwJZM8qKKKgcpyEDwlrOEfmMZPFgM2ip/
gtu4flGA1nMj6BppesB+5shLtaFjNNFf1FcAdf1kJCIWS1N88y3OfgzZuC9V94I8mlKT3G5zyoGi
0xAB4ZkvUcUanudRaJqv8rSC+gltej/2Nkw2QAgiwYcskjK52JsKkGg4sa4193hZVbdCB/G91xpA
jmhpgoUk4lo3xhESAKDLaXYOfw9EQ+95lCBbfcxYBPviss7ou0swLy9oXHROPBzYwDmkEn8d8nKh
/DkxV4x+L3ILM6I6GjNyY77ImwqkehNk1DsbdQHRiOILAgUfcr54ArnmMspSRKDn5Ah0gwFggOe6
8gZs8KQY8Kc1sSUOBzK4snUijp9Ukf8slvik/3tYxDwjJxeIA5ebZJ2ff0j5motBt3dCdSJ0DaoY
uJMa3ECES3SdbrNXlPHB6lcsPrJoQLBojosDWogAXZwUpYP+A43uauJJBt8vz4W85fUD8t7ykOCS
8y9e8pZi7PWF4sjuajDAEj/+xzme7yZvFCJ8R6la/FbruaJ+FLSuIU9z9e/IHnFpFJDIrxfniCwW
LKd0gaz45RUMfL8k5cmcBX2/ldHsnF+sS128KIxAOPtXWh6Oi8WSxe/bTnPoOM/4bJE7kReWqB3j
So9W9I0DNUYlR17yTrB+zbKUUPMff5Y6VL6R980EkmibaJc4COlJHjs6uQuMvknLRozYf67DSDDd
8A09bvKRuBokRiwEpApN5BJsjmW1mJXEee8E2tXWGDMMnVrqsWb5ROKDWby2jKi5BdWR5+F149Tt
+bk160nZiHbz8sQHNtaEiUaRn7uKx2NxJQrZsVw2kjcAif/Hos2UyHwU/+G/yRCjfIJwFrNCzHV7
ifs3bzwS+5WR6Mv3M+nh5yCU4408Z8qUv41P7MSmp0U20+UhcR4RUGr4Xn2l9OXMHJDyFvNo6h2o
8lhlyMJOFhb0iq2GeQ/A969DNfVgGhyCsjVBxbxoCWxqcEN/s3VO2foOcOJMbqeRXFbfSVfo42H6
lMT7+uYvRPAwhpA66K42TLgVzJ1AwXU9DRwDhcpSxxOS2/dghRlVDfERt0MMb5JNFAJo/XSQwLh7
wVeowR+rOBHIcgMGktMwnASFaSmVPL6ffWLlYtVKWhwlUXg/WDgEcH0RVLpZnL1fI/szQDGtPoWu
HpoMDWguppQhkHFe4tAA+hvPCKVi01XLeYO8hwCwYj33L3dymyyoDUWqPJ71flIiSgMxy/tOqdAx
i39YNho4JHcj6TNtge2nRc5ukHoCKQ+Q/UKhLWmswVoTXGxn/OkAVLLm0GBq/vQCH4WqlFhMh0hr
xofdNXyaKOW1Su64nl093Zg9crQqtmf/b9HAIBnaAYhT6xPXUwOh7Fd6YoAqKtdNlkxz2qUuBKSO
uOgMUEYM8MT066O1JAkqz++0Zscw/cc5WGFpvdP+ik10GgL/4kEXSw65eGRKL1pd8eEZaY1+b9zS
FFUFCBIgQnfIzuXD5IkQ/K+GGHrP4r4AJJWh8mdaEnqRbWoGhMhjfM5xVMJKlvn1G4813BtKDjgi
TYtQ5Gv9NxyYeBVaK9+cJlFh3VRCZ3jEz1Gq+TaR3zA6Ku882WuuAElq/LmiA9KO44RCiVIM09Jf
pVlUtSs5b/4ANc9SyPlp1fegFb48uHWLBVz0DmferPf4lIPYKzvrKWr5VIaHzzldS1EBnYuIjmSI
Sz31NIuvnR0pcTD0SXWknvAuITsCBN1jgA+Xjx7IQ3Y1aK1IViuPJ5MDTVKCW4rzIIMdgsDNvl4L
g/EkdR3kB2nO8AG1MNH88brQDUE79OpcU1hew8WVaUI7sHoxWqHrI48spn5c3Q8I4hNZDdi+oVgz
ouk3fKpleM49P+c14U1jU7rXTOR20TEl0BXzUpvQxb4iB1Ch+bWBL+BzmuVmT5X4g0dV08khHVUd
8XSjSPVbrEaLQvbCMGN3dbC4zr1GWIKWJaS792XihMDa4k+42wFl7A0ZbBtCkp3Nh96XdhzQen/4
EFK7TC8mOktgvk9LIhx4OyPDEXgTYf4zIkB3ueWL9I33DOOkEtd9BdDfExUohdKtXsR8m/NkGlRM
1Uxa9gHBq8dU19tXVlVLVLFwZ9YgeZn9QRTNvvWTIZTfdrHCLCnBIs33IDqkUEBDEC5izFti+rjc
4rYqbbdVn1GFUH3aji76ZlQ6GdehBny9+GX3aV+opJh9tmjG2jPFkEfJ06hwQZDWfIUUupvDJj2S
GtS+J0LreRcCzUDYVfNKcYLV138pkXFbFLhPBgBYPgeBeyK+dyqxb84J8j4E/Fgs6q0DMYEbxUxZ
4Muj9vZ3jUiQTC7J6RsWJyQ1xpy6CTmy1qllT+ZLSTiaCFELdpvjthhO5t1EP0RVi2jqIeyLxye7
BtHN/kSS0+HPNg5GgePoHhn73S+mUdyj2AWuCQvsSK1udUpYwgX7eSzgQi1464juMU3ww3S7+mjx
p77MQTyKjKfgI4TV1rFb+uL5SZZwITuMxfhDK2Svxxb5pDQVQOMAhsuUgguLDfJSAUfQ94+IsV8k
OCV8eTXCvK1nsNBbB1O/3tZX0Fsrc0pBldUourEJD8V/T4e8prAexu7Y3Y37fwj7QxvC51N+VfQL
xYmpZpsGcBk/AVSEK5nHkHBPjwSW/mL22pEOYJNaX4CuDOgiH08knbAGuqQd6/omBiaPZWyg15y4
G60skMuBHCqkFmQwW6SRZrNqShGf6OHFELbSsoIYOlLXHLbvtWDDr/jTaE8JKT9mWI5K97XyzsRW
OURw0ghjOdC91sifm3S1dq4HcZQ8VD7dYvHjipGwBFy+7demGxwCFsWKdZ5iw5RaW4OMD6q8VPBX
hNuyWZ1ZLvhN5hk5o26ycnDVk4ZzqdE42knQyI/D7/LsZPvJ9+JjncLH81+v7kheJUmtHvgntZiN
3/SeiLR7y4xjr5lQoMB50TcC4WyGW93ziBjAT1c0ncGrkoYNMcfEqbGh1ZRHarhPRjcOHPZBSu4F
bqQ/BxMouXmtsMZu4yuIj8L+cPNDpsoJLPatnMkIH7Vc9SdxRmvvmx10EYVotPSmWXaMHgS3fDqG
ireWgQ4t6vAtEbiGyrTcXHMoXA3BcHX4kizyKrodzkEdeoVRQy/zVHR6iJTeWaD7SXtfq7103JTy
a8u+Mjq2PQVqEl7jL338RR8roPjuqWOdAsl/W82osxWREnHjl0jpoHXZV7Obx8fFdmTcQKdZPxMN
iqyCAU5Qap7XRoU7nGapi7/7dOtpab+/nlZxBKl2mROHeGqU301d5roBufSzCiyz9SpVJD1pfTvP
Mv2yj68tc4i4b0UD/dpJidRo5IQtoqehlCsRoQ4wMnI0rXfUCsr9w7ncrdVKn/s5X44BUodiKoOx
ubS02YihIGNd46jnwCxDNI8+uacCD1BTAqW/vn97e7hAkRem9uhtRxRCRLJlb3m/cAm2BDOgGTVG
DYud8wCCffyz7ugHIRX67fSgWi3hhwolO+cSpoUANi96JPTxZqkX++K5AFVlH4H+OR3O1TMPS9la
w57BoI71MiUdT/cwSRZ9WKZkr36glv1fBzcj3JUnsRELUkrcQk/BHVq+bs8WLER714gs/+rQI6p1
9o7cbrE2TBWolsLehO2yYVXUQ7uRVoTYYBryxv6z0hMkkquLkg2fieDT5hcL1F7PeMpTlv9xOXAS
PmfHZsPSgTv7TRMbRLLrOMXCxWxiVryYTJ8dPseJ0jKY7YDRSCPDSiRFatJ4NBf1a/uQP75LukFX
N/nVXiJqg5VQqDpf7jla6+kxrnQilWzqUMuMsMPPJFWNbIKNw3kMIlz/JzH50F3vHDHFwJVn+z4+
tvdUzwR8DlMwXgPWxEC4IWxOg7kxIoFGx5dKgQssbTqrwrCjC88IoN3loS9Me0KdUkK9dN4Hgj3H
dsEh0MDDUOpY/oMGy2bpPSz/BdDM4ElDhyHeetOcY3Q09jPgIkLxHVQtdX3neVNun+9IIDXzTW+D
ikgm8RSeP6yWIVlKGAR/pBXEvoi//0oSkNAw4t0wfvGU/1a+3duSjuaU7FDVU6FaLBj+GGqN8VtF
XmI3C2v7hZmXOdJzcDTLpw54nAl0kRF/SO7sg7BAWB3C3/W6yBdOUcMWa8Tg1INnu+Z9qiPd49Qn
oQKGt8jdpRXdtgMsPnquN6F+/9hHqtHSXQOu+91f0MWT5kCGVBY2tH4oIJvOvOLjY87gPd3TaGQS
tF6AIrk9qRCD1AMTn8goenSJFdN3zyAQhuHw/CAo6BgrO77f03uhEjMnYPzJCxWnq9sgVOvJjaWE
eG9CBbe4jcLFkEVg9leWratvalnLFe2wGVoigZAIbxhx8FITPvimnFvZElx2xCfw8yKmL2YBJWLm
h1H41ayacnoWXhmg2x9dx/mC5Xk3YbfNvv2jOe/Zwf9zi7oMNRRGo+Pthjg4qCYJ+WzibQ5QFzyC
kdCRxeVCoezK1Q/cSe0Pn2AzGoAycdobGawW2PsQje0d2JrjaqO0St3rGtrDmOPDr+/+DIriKU0N
xFQ/K7308xDXzSUIzWPBthjWpwF4rnHnW0hKavBJyZZE3Qt0GmXG/JMG6F8kYHqM7ApHzMBXH+/U
mBOPQUz+HYUbAZURd+j4DKLKp8QbXtFthq0YN17KwWpq4oTnuKcHFBhH77XxSHG2EogxyxHRArhG
HlkRuWQOFtlCdIU0trw5KjHt6yt3z1iN4knRV0hagK1oojuOA97kwT9+6D7qTKC1vQGaor5axl7X
OfQfqkoj0H3gsAKMJRl6+wYMhyZ8NH0/T122QtbPDApeyUGbIHSMlR6ISd6fDQLg0aszH+FMdm+j
rYLkdCdPZWN/aKCzWPV62Y06IQvaFkCBQKS5dzO6TUeAVtWZSomJGZGEnOg6KP6OuwK+n0A0c0zV
U1GlZPo850ip1pjNGAhQ5xuT9tHpUbSaHZN6g2b8as5RW58UYhx+zNo4B1gt7QNbiYqU2EcwVSa2
Wj1E5FO65wlVvRcnyYRCoFfxFYXwQZfRoT9xA3SUTo/a2Qlubg96J6pueO+5pNAPmz1QDswxYM7F
K5pQEDdbTVUJhRhHvVdZnANcVi7UoYf3ETVgaUlm2+IRKnd1YcQgyYB5aOaFhGfY71VhoqBeUL+6
I0RucD3ykrLWO2esDLPwH+kWG2L7l4QfTxuTwaaZrnvpTS67M72qsAjaNZ+PNAL4ToWeOYOh/dy3
InPYZcDkBdEyfak5q2PWUzcVLDLV5sO5Y2Qn9H09Ipm5XoVWdwn9rXHOpqfeHzxG8bAuTRIovR6W
ntjbSebMGiTwwbgDomU2+opXoKMKzGFVIZ7G+U+CIdcJ+FhpyP/sfaaIK9tnppxDliJcOxGdb1CR
U3/u7ZfdmSyVFX3N+8krRr/o3Ui+Cci85NJ9m9Xll3zrKsMwH8T6/2pAqu3qPYlCSKQwd2PBDTg5
JFN1OMjCwQm83bg6YhmVnc29uRt5wUlxpop713Y+FIMimSD/uxhkVBLOIZS0mNTgLD/AbWGL638f
w5DkskaKrEG0M6Z3k+GqANXa4OhJtsvAcyDUZnzPzb3HCJ5R7cEk6cdN4BxsV1xg3rZIZJIxvhCP
wxVTIT2eiZtvFa5rmiTOM14QRjKr+HqCvJAR55dR0AndCf/WlU9ytt1VShkmUaNPeIArEkCCWunA
qs2ePm243WXaGu11wCcvqvc/QTpIa2rSkPwpufVDtfA1aUzjTuQ+ACAxIOCuGwt4ahw/m5sqxcOC
W565w+0rT1jJ2WnWzYBebtyNDFHnb7wOKmy7ZltzQyYx1Vm69C4LWHufsAPj2enlgNWy7ENYZdUx
s6fxIMQXbWy4CgXpgWyamiBn4+zHUHG74a9CWwrsCA/DDpgcBgfGt/w9E4zZko9BcFeTNVJg0p3R
bW2D8l36ugaVrzXfwZBzIM+QCvFlEkeeXQjNJBXTCaW0pscyHUtSAK8zlGHcLpVZj4L3yd9jxAKG
HXLosQS7BTRzBWb4IbWTwirkpGOEtCU5buEERTxBdbJDLztkm+1oWpa4/VcM9tUAvJjCzt/jmXZW
HnZveLreNe354n0fBDY4Nm/pj/QMhQPphYjFrr8zvz62AsZ9o3UXv/7t+/nGQh1fTC05VReQjk7o
XqZLwEgLolJAXs1cdAeY+dF6rfWtybap7eO6a5lhXU31a7/nvm0pj7ZZXOXWPPlzYk5QTXbN1pju
xXomHaft03tPF/wd9QMcLT2ZMwApIp34ch/ZmugLBS5aUvJmuUbyBu2SDh6ObYZcsqPHu9R4Dmjq
Xvy/v7ZuJvHNK/mj/8vocEoFRrW2EFUBJ2MqCDFopfNyFRzYk8K5ucLKlbcZQ7KRcbKUWJGbQCPa
XaqYv34SJcFMTxkJKWnJdIBKKXmQX6NVdDeIlVXKwxXoMlH+hFbvUphV9hXR6b+S6+NBQ5AO8z9/
pEB8XZq0CcVGr9v7zBk3wAjdNBrgGbW54S4KJaFf3xlhOrn1PIBAGLJzhBas64XPxDHOuRg+9RmR
oOs+rIb7jwb4+GcDiJ0CdSqm4G4/1qkKrIRAJTfFjuIqnt0rQyOhEyDAnIN1s4mQJ6abA6ex5rvj
s1b2oIpW68gFhEErJq9rsFqn74k0Vfnf6mI+Uw6t7A7PbPhwWeBkm4OTCktiOeoeamTeh8Udske5
cQwOV0OGmCv09vOCZ6dZEwQYODTlKaM5V1Qsi9x6RI6UskA1SwuLQVT66eIfNmGxxml7wDO1aD7Z
j3RWwCq9Nev1eQBy5iZ280Db5SLLtNMx55cq7TvbJxSkdbIrvCPGmMOWwegh4oIWOpy0vB7n7c6f
WqzSAPzbFwrcbpYGQS1J3v3uD3dI1z5BD4C9Oo3UvtlxH8JqzppcRvvQeN1VrrN7MFqP04yEdygL
XKizxISbaAoQTx+Qs7tMMQGuQBvsyff4q+tFvKsaj9B609Fh6HCKJKHOm6E17tNAgR169UXKlmm3
aXo2U2EhlB95qgUFSSQiNWJOkVxM2ASGwtpOJLU1hjGwCfhd0yd/oQmbHiiMMxzcooLLb2Lef/96
+h9U8fdkZEsmCDANlToB/GPkYzxiWGtqL8+60gfx/XYDAuNZOJnYHv6pH0aLB58zBMo3OWcG1T85
xEnNMSbYC33KuiOqog4aweQFGBlG1qgMT8XPmXIhHH0tzpZMTDkzTFyYFzG8/wwvwEY5xGAetqTg
+HxYIVaNMcTmJC34SV23WHhpScvMGYwt27y5nFR8DTC0Sa2Qyj7Ho+b/mkQ6rNhmTU/DPLnqSb7u
waAW7Qe1dSy6/4IRxgOskGkOOwYbdkS/bZ2yIcish07Ae6eVHemCwv0nll5tFLx5eiWV+MGgO/71
7r09lSf5xT/eJ98sBOrbXlXkzueOu981t/cWBJEKY4u71d2BelZ0DSIZKJy8hHBSMpZCtIDfYYDc
1GCWxwS8650BiMhUjH1qwNVlMJnh/qAz7nDmKAb1ttj7aUWrP2JWWkTieBhYRInZzI8Pm4TMRSbq
EWK8G8uF1HaWIM4k/gxMbH2lofbMBhWAcXHJ+Zh7NfZqMdwLE3TI7w6KMZHXAV/XP90GFtRQ04E8
BHTaF4VPrLBqdM2G5QIt4/AVB80VQmralA1JJbI5nxZIojgJiUUwZmSnTZtXB2hrK15KF1UKI0gl
k7hUBKAnVhPMwQx4X7+hmcNXu9byX3RMAHounw3fMD7uvWwzj/P84w251sY+7BN7ktbVI9f6NI+5
6nxH63BuQ6P8M0WoArDOYdfgSKkYQ+0BCHUoXSaj/wQvU37FmVTS4RbxiHCNH2N52gQIbTS7K20x
Br/gxY3czjU07oTD9Uv31WYRspmI7mBj/PMpQd57H3y2eV+o0K/W+aPVzkgr9oXoBA58XHXgRJts
c54/W5XWxMkywxHw+pInA04AM6Qq1R8cm2GQlzCKzKMQ+7ATF8hpnWcnAYTMGK5bM3O1r8pvxU+h
oaMvKsjGA8BCpwSlfmWpTRrtH4mBiQJrl9dPZlAIBwABhc/j1PmF964Ub4P6YTVFDcabqjAoGayV
ZF7Z0gs8sycv5bRRk9XJetmLoDNnjpU4MXvH+LN+tc0re8RUMs/q7fBtOLMotT6jLT2fMa3Ca1Yj
ifGEYhwvkm8kU64P3b5/5Db6PD44Fgfqn9LQp5FOR5puMZcGKoD0KtaxRW0691loYMEyOIDhQ9FX
WD//VfMYHo7yl4gupI7FsNkOjjiIbHC9w2ax3CID3deNc3czvLNKX18Yuq+RU1LeaHDeW0D7tXrx
DZjnZA8jgr2wY/Po8gSo/tB4Uzw74U5Nb0WQ1FyIoKgBe0aLhAAlHcMsPIqcYfSnjzj6ML5sXZog
eMEOBtoXmjaVFZ2+2X6zDF8sDfmFmIV31WJCD7lBSIXOwh+4bujq8+5qLz7ZI5mI/z2SMTxnvUk8
6zFD+MTHf2MtcUqQwWthEIuzsGfGPD85DSQkjVS2RMXmAj532UyK63kpCB6KNB6ZRI3Izu4fugz2
bIO2XetFiNJOOBIYi3ZRRwszqCghUKTb/Jd1jsvLnbe4mC9TOr1VRu79RgN/UX1LEifKHux5Qbhx
XJ49C+2E6oIwzsU2fpGnq9EujhQ+dY4htNS2diRpPefCkoInKvLKSid7d5iPJjPuj4RnUiDW7pm/
/U7hfv5krBCm8jh9gVHH0Dbm7xAWpW2b/TP4eoqrQKprcdL9DBe9lQG1qROgSGWDZ/hYZsmVBBWy
E0XsajINE50C8qV7nOGWhKE2RiNZHPQPzJek5m1+bAv5fZuYCVZBONNzfhtrZnff8acdQAo2H7EC
qdEfbJn4iHlJoEa6Zxsfd7Zx7TG5wD/o5phzO8tMUWVyWyDz9Idbtmf4ZpGs5Yav777dN7mAvVBT
iqG7PyHAqtaMMO8lRnYLBW/SRY6NJeXm+KjBd8uO5z/uSU+GGS+WWQvA7Wtb6TsQFvYkNDngaBdW
kE8RRIWfy4mUYXHVuFuqjRuF6xjaqAHC44eJwN2QsTgAmZvLxOl/e0MMNIkYcaR13cMCwGFqZH8w
Gwp4K7C78/ni8xRPbOfYaoupo41Cy1iM6EoieieNrMR9J1wykXyxE1Rc1e3LU58vXS19WPWpvdeq
+AVerXTnqOkSlAqOEq490UNamM5X8Eg151vZTID+e/Vq11oTruFMibnV1xH0DtqZ2ffouGjbaQ7A
AF94vDxRGT4h/J8YB/kGD05U8+VakAsqSb3Ll2iNHA1CCimVLt/4lM9y2/5JFV67FDaeXbJ9IiFC
RQp2d7WFS/E1dyHo7x2DlVsAn6zPu660Zy1wVscDHfpYB91ndi7N5O9ilYiqLiEwq6Mqz6y91SsG
VwaaKwDoA5fuQcrV4zTJRVOUYb5NGKH0rxxLYx/N36eDlZwBoeIBnD4VSrfn8JbeXFDLEaUmYwec
VfPPRwepVrVhUhRWvrCFPUpue3AjKG9b50xgBd6Zrymzflh/NrwGdcvZZC8lK2FXBHPtlk//+VV8
NEFM+HGWsTFRdOk/QTQ+cgi719o3TnCKJEUIX0HFua0PuZOik3DlxJQzDbOVsrumoz8VoC6NvWGx
HJqtloHvTkQmaFr5hGhTSbA/snxnf2AG8j2sdeZV/Yyo1t0vIIOISON2FaQRsvbDE2Y7Q9OLs4QW
msO3wm4Yc4sEE+t3iq6/JlQ3IjkGq3o04jmEsbDUPy4UO9Ombo89JytNzYir2EWXAHU/zbLJu9Xw
PVrovfExHJxyb/0xO0pJCP6rlLsZtjd7WvGS/cQx5YgxrdF6k4s13gPgvm37Mo8Vs8BCi2ccYFaj
h3Pag4Uvxd7yE+NIX3bKEgOrxyWJo7TrmmmhE/+lgdRfiQEHQZHpMmY9cT+rr+W5mDcPEGnJYXIr
/GexSljTtN+5FzPNRYgYmfnvvKB46NZejO3rnAO4Q1SL54CAK9oJo/1ZgTyz64phvSpahSxxQ61I
1misGMc0E22okReJ/1xQlAY2Oi1t0zPDLFnkYQ4OgpYA1t30vXxZgrd/9dHm6oWLRA9EkPxErntn
JEjKEm3YrsbVe/d5Dg4X3g/rVKl7+9r3oVgoobx/mfoXM4tJgYEILDwZ6aMGNtErNz0dwqcOMJHP
4GR8jCfwil3LSE9ui0wzrpLmes8xvyRYU96jC6NYAUhGbET1MwTUMoIObLPaSTeVD2Q2KE/L3Hmp
C14aqYHKnCTxW0IeMGtJLyhof383l1gGNKNP0eebV6kVJsA+rr/715TmKUQW6+nADmw6ImuXWh4T
S48l8czhCB82yBpUu/CjtDQmZDA2ooH3skdqPUvn/TMmwnYN/hX9jKMIM2hCF2ED8pxaUeWDpM/i
Mz10YgTVIm5nP1LNYN4jTCml/0cxSh3+sQPSW5zdneKoLLFuAbOnyqt07v8rGijVG/7PooZhs3Mv
bpslxtUC8TnIpJr347oBOZ0/FRMBjcfzKib+3xmUp6xp/BlmLbR38+J2OPIzOm92gZFY6473uM+c
UdsFQtU0fi+YlTpuI04Ngh8jmElO4ARPPcbzS/rQsUPnF86DFOWmXDGU8MHn0n58ME96VBeFlipW
aHJCaMwGKdhq8BAANN15CzXdqc+36zKX7AqhW0KvMnyg0E8CYb0Qf/Tg26Oi+ec8+hGQ4A8FrL0N
/qvROxVs/gZFivyVxlW7h6pIsonlRdjkq0p/cgZLdq8kAVGYQ7dqN+rXPc3iLIZaPGHD6eYCA3VA
AWzRS+Fj4dr+3Bb4QygB2D1j5IiaP8IWbbSkMewyXtp4yKQ0nUuqo+9YweUSHl9LI6cBnt19XgxV
Wvtcg9GAT8tIHocVzdwrywCFD9D/7sPNUFZVjkIMk7qQ7Jp4dY5x+4YHIPLZhDA4gJEVqL6xembY
2VQLVei5Q7LU6xkdy5UCkA/m6lnaIqcXvMcbkYvN+nPSyFsk12qSyo2siE5SxlebbAl5qNzRdJsq
qB7u5YjsHOKE1Qs5X2m0iPtvE79wSo11zpx2ZYo+gDXJnyoEdYx2R6cHM3b2VVtZELDWvPnpqDoB
8OsmXuZ3kk134sLkWXnTLzRIWtUIQe/cMfMkSuZtC86mdXI2Svp46+rOFACj0ylqET/lcT5nCcbV
MX2igzJmD9+D9ZUbKYNfrnGzdZg0t+s36rvUaEw6UWTEqOe2qSIa91QtQusygyXGQ8DLLioJ9O2/
/pp5dOFXMOP5KW4AYpk9FmfeaU9mR808eH7TFW9NAXua7Hc1K0rn2N9auZNVr2jnGMsz2f32R275
eBJblbDNX1ciWIwuwFzcrNMNlNXjIZzP1MbyvedztYr0jKLx0efQFLTJxIqV57WiMVzY7k6HZHcr
vuT67knLIZajHJhxsMLLIcn3XdNMi3PFQA6IWj1juI+X3O4feB7JuYVUpL7Na8h32/Nd3PwPk60v
Nomoi/pNViqrtXJiHZHBdHktIt8UMa8z4XfTZF/9FCjeQ7348xN2L0uMqKmaY57mks+4Ya07WvQB
9465vyihmErujdrPBceAfpKqvMTy3pCa0tbAAhLFWQu4Z9vP7zbz7vJXziM2gbprMyunxE5zD/qF
ZK40MHmbwzFe6N1Sb56PH4QeXGSOEnypQhnqzl/4Zljx0XVd9X357l/J1mWf5pq/D+qksyC9KxGU
u/FU1jp2OZNKD1W8Zl5ZjJHP3CrJWZnlaPkkE590nEZ9YfUb9iQ1WGppeQciHJwcBNucrAQkUMYv
Tch1mRYp23OCKQcNf+cxhuuQpyZW/ncfTi+HWeJ+OloD9TkaprAixwlB2KXuUCB7Yuo8j9FOSDvx
sgT+VXAsxtFJf6oKWpN2LVTh5OWgaabMRA7lvutmSJV9t/V/qT3K0DCRV5L2K4m9GDZ1WxwpV3KQ
k6Z0pdjLOpRgdKCNeYTydawydTy6x2PvLIbMJpUCwGUxqvMm3SWU3PKCVX643AFgHH7zg+KmIq2V
tukx2tNHkfyM8WYNjUsp1rdUj5ySe5t6KIeBOgMT1SAhC2kBryL0oo5mGbiyMED9qGMJm38dkg6K
x4BVShNuSTLx5i4b5wAXH57xINNgRfDXSiKLfEGF78KDrklQuSW/CzIpG2k3JlZ8aUTb6v/KKjzy
+PFAq/Xi3HyM9cGAe+dVJ7zBBdXimBs9qhUOJSMh37TVzV7fSC7qtwqmCHRR4wH5sfbOkyNNIrCC
wYjjiUNNC3p9aYKxXYJAPTD6ZJCQ8SjQ8yBiQZ8spaiV2KLykPUbRm2HaYH8+4e/GMAiaPjMLuEI
5ljA7NgnFanGetK6+nEF15UheOFGGg0xMuUKZdqotT4l6sRhpp/ccnUHg2s8Njn8h1PIYiUe9Hk+
b7NAXdLivGuoPRWJ0AdEPnkRZ4oibKtPXg5JaYC2fLP5+Hk3bIYEU5yjCxee9TXFrDmNfa2485T1
v8A+5M6m7S2agUSMRTmX6TnGvTLiEev8r+2Bg7hSV3pBs47G8uZ+YeRI8k6rfcdu8VPMnTwpOfAs
3+8a9HnqIB1W/okm6dRY10gMZlB4xW+9P0tZrNjmU7V1L/rCoj8PBpqqwJ3pk2JIDq1I+Smy1e2I
eVjFSCETGGPv76zHDjSaOtgJpYxtJsXbceWMVNedAx1+BP3UUmnbHKg8PLRedD1f2felPSbdlqTr
uet+TNn2VEX+ghJPGEvQGD+LJ77MlEV0ljOudDcgUvgUBj9H28PWGMbvaBd/r1jQIEl5TlkK9jUS
iG4T8XxwUVPVV/UZ9+EGM3QkIxASdwgj2LYKrqFxVhLN/2YEAasM8dQSD66AZ4ekNBIVNvBYrgwR
YFuECeqvSOAtYW5IX2P0bKf8STJLz05albYxVVn9++rnfw0+8Ts6snf97dNAwQ/ITeoZ8mawalFR
55s5t+6IgicZAx91oGSPupqBH24rO7T2U8Y6wAD8Iw7r3+pVoJQecZNvxXWI5XVkU4+aNIqKRDux
ELNt9wgZSA5UeAXH3omGnNqSpjrCv2aPZvsXSaHf+d6vYA2+dAz7co16cd+z7GNOFR9i20iR3W9G
dIzRz/HycWS7bYE7zvDk0CyXqvUM033MNW7Mu4WGgJEN4fxI1zmr4GlxdRs2c38aD4NdhVxNu9eS
smMriJkwRPGrV/ERw7kFPFsDYe+xAQhp76TIKRsR6L2qdLxoijW10Ik2HKGR+eyGONUwxSJ1ebb2
V3YhBXGNqGMqTBjX1etAuWakjwfl1FubYAUuFNvABbopFxYhzHi/TMpcRWmN2iie+7E4qoo3e/bp
yP1KF7iz2Aijuj9KWSC1t504UrCw3uPGCcUirdGVG4R9EvbtvKDXV6ZVeScScZszr1u87RujUETI
Y401QThOPZXf4ZiexZxdbQUmAFzJEsXqNzrfTuSyoMfsm6lvdOIPWiwmt1ZtMPYcVGMeRbPE5fhJ
5F38lHeIpDzpi6qhCN+tSGJO+U8q+r6cLMcDUkdJ1zfjLdFQa0PqBCkibrRyln9Ia44WPozrqFAN
P5fDiqPTfm/AAFLQAQC3hns3SRE8Q+Xf3eAomZ2HNB6LCRefcODRTuGYv6EMYXAnyMWw/SQXzWtD
fWIfhSKbugGW5SwURg0sGgARwHiiRFQq/TjpW0VMI1ZNr38E3k6NrVf1YovaWvXfTt0tK6LB6Er9
QwbuVlW6hXuxBRzTohxTj2WF/CZ3jDWGDfSY+zCYmlGz3gTiCq3WiPUVzto9TuO8QQ0iN73M9rwN
Hx+iBFbBIqH0I5DDgid8H+gfGS6+oXrTwdTXP3McswO2QdEp8UL9kYA1E73Rz6TzxKZeb5KVNv1H
Lzt7fMt4GPsl2TtegbvXji/GEmo4w4VSy9JTmF+xjbt2pKJARcGp2o6yVLNT4o+kDZ8pjF56ksTl
NKXGjdUQ2g6PCV5fdkVRQh0T8E5SnWPu+hmNkKvsWUMUAIOlwXuXhvvC6XQbxtrtEg8DBdBEd+7z
t4vJ3fCuAxxzMN6xxKg5PdM+Gr+azNtELWYYSU8OtXw4VfhMuGy81BD2tb82l1s2lPfVZMig5mwQ
W2O67SYo8lXS4zYIf6Hb47xTL9FHLoTmkw60IVi0haVLCfii8zUdWfTwxqmgd+N0nKaB5L2xWKQT
FNGyW4IRT5Jlsz1pHeV+muuEcwdZaVzXU+RSij6jiNRE5TKQDoU74FSKD8pf/zm1NGY5Lj38GCfr
ILiATWqLiiZI495eKGdAY6YUzCpMKn0sXJd7spmuHajRdWslVxE/aWEU9kDrCiIXSjqWTFmE+GIG
eZj7bfa2oaQAjFazSCWkpseSyw3TXB5vnzSSBgPjleRyTsfLmbFUWnN+lDpIuJXSNBm3ZBYg5RL5
15ooyzhBw+SnqaI6m4itN9JT2Z+O35A9N9BOi0jAwtxVUAEo53xxLTwREiIsinoGdpikAlv86+Bu
27mfwNSxyqPoVwaLh7uvpgRun1t8rIWMXFZKZQ5d9N1OO5RZb763sxQt2wBeU+LiHB7MfK8Kxvlr
yOxy1OfnaHD8Q+hekEMhmT9pSvjzuMhqJtPU48ZJtyN2QqAxwL7G6FR+c7rjhWZ4Te1TehjT4jVO
uP98CeZm+cH1Qqqf/3QjRdQI6yw79b4bddTfVmZ/cTiaHj/dM/Gx1vmJ9HFDJEIDWQPfMn1P3f7m
+WKwP7EL35OQSUq1iiHQR3CLFxzC/LF2vXCHiKMoG1ee+Z+g50Vlmf/3Wmj17+wNGeP9r1sMGP1m
Ij4vy+lscLoe2Ck1SA8uRp1U76syJ3Av2iMDLyfL3xOaIbvRar9t14xg66HI7mN0T1z7yhn/zmaW
rx/DQJt5lRR64Ly4t/I2jKc+cXUZeco2M5yFJuZkZUjabZcESOu20cS26qE5rKItp8w0Y6SLd/9Y
5HQ+0qpNoggJeAfjEyW9xgrc7ftHbkUBzHzwoX5lDD4Pv+vv9w6M99F+IojdyUTUcRfqsLMhejCJ
5qCz9jHL1klx8OxjBSMfgadbdHJdx8bJ1RCbXAQey/U2dF7XGqqsG4WavF/hyPLbg3AChL9E0hxx
ZjfpTk+uDK1oFU0j8AJ9xnfCTYMq3AbROoIigSTzqku6FcP+IkMr5soC6IlYpKq9UiTUhWeop/8v
GnuVE+m33qVCVYaMMdYcQRRGCa94E6tGR2cfEJACy4sSnCHMAqn4LRpMU2JxeCdo990nbYRf1y/P
iJD7EJr8cK4cHfdKEkA9EXWgOfTSXD1wuuvk/a4MX9Ok+AwzOF8KR+zPM+oO7TJFZxh0U7gyR5KL
wqJMfaOiC6n1f8jhbIac4WntZRJjh8CqR6WK6OOK6usZRBsQijoO+BOs0zTQ9wJm+6mjkz4FDBDT
lu0RtgVw+E3DCG8A6alc9eVMbGuG75zBAoE/dwI7B9gzT1c+sLFpMrqVhJ1YaYT5jpRdSi7MWT4n
rv9pqRdLswku9rthUrFTcqlkdmspGHO+/thRTqMn43eukaxmwjkGhOR4ZHPlmIVlbnUFexZr9mrn
ILj1cf8RQWHKioKvpg2nn+0pqKeKeeTg8Wm7peVz45PHsss429IRBwTF733fXqX40JchD8dleFBE
WGuQqsXTz8z8elFQYqmRmjKGH5j9lk/QjMysBkF8mHrBJ6t0T9YmD+zGVKbZRH6bPBS3PuuVKj8S
Vd0wN9/7j1VBmZPCTHmXIaBHm4STXAYAX9svqrJRUcl7L4vlJ45v7N/Zvaf7gJCblhG23b71+vL/
ktA0ZAAxQs2/qAlVLRLeXs4CEXlwaYYGdqyR3a4bZhrYEnLn6DL9NErQ6/HO5jjcZOYzZMIhYGb0
eKt54Q7vL6zejOc6jWUYKiymXjRAyMpoNjzd2vtDTYsxu2K1Cn3fI4/Gt6aP+b1brXTUHuGubxNr
LcZ7bzsSREkTIuHUhd8/7VOIBTPaFvLBzduz50wX4cVuCU9ImSrIggxMmIp3pKVmaiBSU6qArIyj
i2aNbW52wfzVa3QITWIjnQWJGIHoKu/dFhT8nS83LhgZHSuxTz59XrkAv18EOh5i5SOMA3EAtixz
SNcair6aDBIied0ge4dDR+adFfKMTrny+2LlDzTCpsvRgLFhoa39e1We9q7FFzF9TPzo/pgwG7JH
dGO9VG40Usnlqc15P2Uvy/q8y76ClmccPQjWJwnVy8utvJQ/MvhBdJrkXVwt5cDWvmVQ43Xweeui
BTAc71A8ZeyhO7VkyfqAH1IfrZS7pOqWGKSp2ixVhrFOD2VjvhBGShXyUjAx/VuFswkQ518xJSoX
XFqFaj7X6sfj2NeiM+ihedDK5WHCnsWcHT/crqcKleVEZN9MRU9LNLjVBNgQgNkK4xzlOwec8oyO
Y0xtaEk0z/u8OXBZ17GigBRV7fimGWooDvnFUV6Aw0g0NAz879ze3lhMmPVQ/WEqarrX5BFdV6UB
Cmr1JqzRdY2+GQB9/YCqO6fmahFtrmAIUoMQD2lDGyA7NjnoxfZH3qvF8WMGtGVRxDLxpb+E2X+J
dZdLyfyWCflRK3lEK60TEy2OQ3DDBSr9tn4NdFipA0KeKVz3yZUgri3c8JwQaUkP+EB40S7ye1pV
+jCNXdAo2Sl6/HacUYNjiVjQXpBnqfk05fBZYEF1B1yBPP7ObLRN2xexip74yRWCc4JLb3RTwpgw
4Kdn6H5321O8yCtwv/Vh04MclhYrkdR56cn4BGIGcTHiWP9odia0sWeWCAHO38eFwG4PpTQnJXPa
7JNNqPRenSLfal2FkPd+Ua55rD2pQx9lVkv0YDd5HWl8GftpscbRRj9FMjAIPPGmzvbfRJrJybXY
THf74VpyRjQcJYthQMTkZZ642ODpJZyesHdRziLgu5p1m5dP/dLtPdZWmc4jg3t5jiM3dWp3NVJK
q93t2rzBEdNMh9w2jXrE58PSc0CnWrSSNn31ApuZvcZPScnrRrO4bfk7I92rDVJZKuoLcwwhXzX9
YI/BdZcz6I/0CV5C5Il7nDs0O0vv6yKCMkOCd+V9WlHweVrmMP27Tx8k1Kj76U44EHazUZCn05dK
OgH8+7/zWFBIYFlabE8iSsULJE7Wc5UoEtmQzpuSBpT6c7yUHzUg2n17Vfenq8gTh8AUfuhQVP/Y
OYIPiutCQPq+9krSwvQJ2vjER8LE6VoHHqh82Ad7uCpFT9zlgKfT6+WJGq3pAaechOKVDlkVYFSw
cB6A2CY2kvMV6S1ZzxdrGPoPD1TKUOdA2FzSEykvkfKASwdof68NRsKsh4Oo8wTpBdTbjZ/GTL8f
3s6/wUowTMFMFBjKOm5kr39t7uHoVbTirkvi08T+17QA2RMxKohv3ksy1Hrn890ejFZ5+oDYKBFL
PHoqoPq8imawDezMmXeOiswpe28+kySjjC2GacI8Jf1rHg7UFCDvCRcdw8bihRvxWkTvJqi6WqOF
Qo/cMi5HTvXdbG6crXvm0tRD7Wv9xkqMO6WTVUouCSIHFHbdrqkscohJXQjH9J7zMB74KPXCRgRr
17PRNCedGj2CzKIbWRJm1iC+xmSE+qAM3NVpVGULIQqbSF19wif5jz2G/otzhbniPpVHBEx2GsPH
jB2/y/eSHQN2L+0/CIe3LuQgtlTnjoUqKfMF4OUvrwu7zACNsDE4UMh2GaXEL8XypNKPd6gMJ7xU
CTkGloDSlW12ivg6ivLqcMIRay5Ch2oEaumH9d+qHuTJGxUi3nyzccQPGCSMXF40dsUhTPsGoOSZ
lDqhUV63aKsM/D0LiZkF47olpnqNeq4IoYBSGCoVQ4uVh98G0xEAtQSSIurMq7KD+sNh/2fnaIYz
lIBxuZWYX6iAEPr5IRaR97DEgiCxk7PySuPFPzDkoezmZv4VGfseMbg0a6YOC6YU13BvcGjFzKEd
AP5uO/YVXhuaJpOI1fK4e2U4T7CQMRur/z5cIQCzAan0jTqvf+4TZRnjEuYWzHQimQ6mYhZyrEjt
0eHg8OID4/WKElgo7XAYJFo7SBI1I59jjKhNMMP5Q1KHHg6j6jpE0GLVw0/Fqj+5X6av3J4qVBjN
sx0/gFWycJW4Ft0Y3CXKU3kxNubMoaxoJsRfccdz/ndLWDwXkQTo8QtLJOWGwaBY8tvXq3/xHUxD
Hr2+plFu8iR6Ptq+n8CIQhHOvrDeYA+2GXoAtTUc0SESxFhHbkkUZ136uRm7faYQFOEOB5sOs0GE
XV4ZBjodlR9OzLAB6TtbdTWAI8ILLtdWfuVFxpNm0+vxcFzUEbdYDjfDy1b+hZ9ZuFR1Vj4xJz+b
SlyltUFrtiVo8j6UdavOh+gpu5S+Jg6JCob/obZRrC6iCT9BXMl/OoslM9rT55+2UyzQ6SruCY7s
ROMz66CV+8OpEXo4KsqcLkmUpoQFvUXW9mck1fL9pZx0ft16OTJBVHkE0W+VKQCZq7nImtDUUnhI
vUJjMmr63is6iy28JNzyFHw+Mu1HfMEGhTy9uIFKqq/GPQesBCVwtbFDo6bDDmn1kWbP4/sylxTk
yeRzqYnNuv1zHpBJsJqr6ldAiJNJiuilBgun8d0dZQCi0QBikrPY4BbHJMcYdEYv4rVHtSYYPvgE
364+x5XeP+zepMnNXst12WDvIEkn7YCcBbU1m/hpDAib9+n6iTwB/4BGyR2WnYCrrhUTY9BImfOE
P2Crc4T4Ce3h+3wkgKUdpO/P80f7/Bb8ts4SBX8rWNYsACZDzAJUBR8+uX+bTs2vbFRpQuW2kzwp
21KSqwfirMcyXHx/L2LHzND6l3IediRTy2zW1u7L17gV/WAxsBM45EkG7zEZWMyiNdHxQ82TuC0U
hRvr8rmfN9Vel8mHHe+m2adaHOIuoSsGFatq1mTSmGO7LUsSXdYUSlC8f/Cu5NcLfCKmyWeR+5Fk
iwRev401frlCsJy5qltGHpa2KBXNa2ws+yhmCZ/PV9YW2me7ehJ6EoX9tu5ImXNEEs2TRD2qNd/V
lz0LcAD6IXyCgLXcP+cv6s17zhSjuKqNfo34MCoQNp+/5bDxBjeBRFLXr7ZLAGbb+8jUq5/3xGhq
9VgzRByXlUp5DCThv1oxTh7d4U1qGtUTpmYkIFcr17kF8RXibgId9et5cjRxjqHzVYQjhcgssoe/
1ySW/VMRRpnY5/U+/d/hBWnu97lPKRxrbSzlXbyxOW61g+VAQZVLdeP2LTraF3B0N/Yft5Wbo0i4
kTvDWf2CEz4DJAT6yL4KJCOSS/a4YqK90I1GAfLfkM/hTueD/TRRmMD4g8BWvZxtfBvAtpVtQvdY
CdOu/3PCHu+Xcx2Wi3CzINmffqjIPKnKy7Z/NeMOe+cQxsKGmZgr50kjjHvUUV5LmN/mkkLYuMRC
rcF4/8rWI8CHBQFnqoe/flWejfQX4O3SYbVbw4kn+qagb/XqQRDhySyXSGmFH0wTaMnUHQ1o9Z5R
bS1miulGvwZknXrSIwqtOzNOrfojRW9//E7YFDQCTS1VXg0oSdhn/teujlDA0ZgqtVVjpt54o3MP
ZCidklQJIClK6L92wesCShKo5IqX2skyKLCdKw28K0/IrXYzjk5spAWll7DU3JE3tX8+BTPE7Cz0
LEBB3Vjd1ROCsnaEEODNed2wGxz6ylqAKGsZUUHNccLcGHntNF1f0yQODRksw57e55Nh1lkc9oKY
pEYYR+vo1XWgRQerIaC4IqvaqMdp2/zQI2XX76NKzoxPTRNtCCU3Skwbc0Tt9aYb0HD+nLpRVaym
QNiHCNZJymW4E3Wnsi3mlUVOrXDqKmWmtx2D2IYjcpbPQZKNqyigSyMjhiwwq3V3dSGOg4SLNDKJ
J1qQ6JYtq/DMDru42Tao04P8pNDCFCPqadJo7nINCBdcBvBzNbLCGSJuZlmMKsQfu7zwCgcCps5P
WHECIzMBnZADeRVw+2dhrlLNOUR0y0sIDcLel58cOwEi1NOaAKn+pCYuMvTUAGwR+Nac+bTo/xVZ
uFvZ2mKMViKut0sm4KHduoFfiADkKfSKuR0wqfzB6VU8GjG36vBTGHvkrgx1L/DuC6H7Z59DE5Bs
Nn3T1/38RCjok8lsZlXQRMl5t0tCYKQQL0QLbLbgX4lJ7TVs+dx3/tB0H/TnJMWbMP/hDfzcX5xW
O3foEu4ZvbivjgicYcD6KIS3Unc8hEy4a012AbEYOaV5QAVyirD3srSKmZ3qJaOAhr9rBFF3gLNX
h9G9ohhzktEziYpgqkKFgSuqPe0iu7M4qz1G50kugCNjovEdwAVfLzADRwKQ3JnturWSF+LCexrS
/TlvR58ggMjqaDr8OXkx+kcst9MKNr/0sl1YHEJpwA899Rd5v9vkuJHR3nEEM3vqfXvMyoWanOFo
btvZRHpVnEAWqg/lV9e7wxJCOe0kTwa9zd2IdCwn0Q1kquckhbv5ZnI2ihVIlcBG9YVceIV0LZ2m
1DwMKzxfyv86WPM2ZESi6nVNg7TbD9IjNp4YMg/QvGcN4i1fRhMwBU9GcjxAHXx1sCl4qAcYDXFg
h1p4yLUIF/0O8o8cGXAGHZUr/hsf9lL+5TA85Ww8e3dYTpoGYYWZp60raWftv73l3EJv0UHoRvpc
cUr7od9y/WvvAzbhSajFgzgUAbM0KJDLCOVzJEchNyV7POLKd8lfcdexvSUNMnMGV1R2GZAhs2NU
U2+qWO7e7GFZovbGjftgKe0XGfnIlUk4ZtAmSY4GOC3r0Uk14Gqm1g+ql+GA6BB4HJX06RgS08K2
eDZbY4E3k6F3pSTW/KdFEQqhNnFXWcqqtbDYSwkPJ9QD3nmtKs/8Wx1GiuOQtXUZ83WdO/JtcXg1
7LN/dNePltmeGYEJe+zTMfiP13a75+5du4vZPzRukGGhAprs0DYbah5zRMvuWFzUgdFdDCHhqLl6
ZoABGVx9sTj462Xh0e9QI00mqVWdbQQ7fJsyJEHD6tMBxfX/jmohGYw4WnHcEmoHNCacKXmvX5Nh
L1WM1rBlYclK85J1pY4wKy6jo0Oj54nChSQ4r7FtgsSWNqN7dRbFB8uzAnxkqAHPEZIoUqDhGbPb
U7xvI2XwKXEWmKoI0Lh8s6e5Ph7h76lTxhUMRKGYR6Jr9Daqx9A2WXXHy95IaO2oFpZp6pnYPUsv
u7Heu9zrORhHLv8XyUidaZ9YQRDI0QNkNzrjDXkAdGD41NDe84PKFPjsBRTFZiONa2BrRh/4Do6S
IP4xyo+P+NO9A7tm7k5h5LW6Ut/n2Wkf6E7vGCgrVh0P2CCQm9xLcsS5ev4wC9ArrgRo3q2p1FOR
8TESSPQCtYNJPi5aDspHiV/o2fcz2kzj5kXVil+LAA2pK3mSBc+jxmIZ5wxTKTMX1kKwumkwvtqk
LAuHuxctPb3coaB/0jtQNvRe9/2JKte27uO5GEnfgn3wDcs9jOF57DhWG8FoDUWkuz+eS4UJLXOv
nOLJCCgpU7K/wXaxXAHZAath1KkQmccIMwResFcf5e7in3EvBnzNBGmNHxGCJL7x1nx3SomZGc5c
Ei0RGAy2qwbnqJ5t4NLrynUK/H6TGGlWKvT7Z9YhMuKjadh+ufVcI+9Fs8JNyoKOFn/OvLkDZgkS
WmJN91oOLoUswyClEn6m5YlXGD3KqjjQzz16vUgtY4Iq5jf4IoqPUV9KQubgG+qtSC0th8/JQpYe
n3r6/INSW+2Bl2k54sOPx+1upBfQhFpv+UuKyhOltIkaVqDuVqQzzPBpK3vbqp5UH8BkVbrKBYKf
zun3lPQ4vfLBQVT/bjpq2AHTTD/0x1iZEPLXClOcwNpeGQPM1PeqpIOqeqy3r5QOIHtWzvyTiCJr
DyrjW7KO7nh4a27qEhyCXwTX9lvcCE014J3I/0vORD3PbYtliKRBZpppuMEJnDLj8K2bOq/vb3TZ
b+U0BNv9SFEMS4EX/JLOROG6mekk7T9DdCv5ZvykkVoz3NSFRWqAAgSLc95KaSAvcaAtHX5hwc7+
teNbP4u1hDroQan7UeCc9d+27jmaOsRthCvnr7V5vnuI8wWKvFXNF/9bObsvFhe7/FILGGt5sWqJ
YrKGz3m8MB8FT9KIPPN/bDj1DiIyzTKsegCvg35Q1sdmm8niUrHGoSsLsIYXvDavp+y4M0oAYOi4
6egF4+2zpyhxjMZDXvaxTHtY9FxGYMazqBziZLWcQclc+/gjO3iMykGrJ7tsFNXDCH55/30gutzD
dzvfQmHkXt1ApHIGNiWA8CJgBs6q18JHnwnFX67a/oI0fbpW0GVSM5m0keKuhwOpLuHSFjkhufPZ
ufFQ65b8Ro4vTs/5UZ9kxqYZidooQfbwLGhbCeYV1ldR5KbHloN29dxnXvQb5nBuAbSQVwypx6cc
UYg1NbeZWtVRmAKRribOktPrV6g6JNfsBaQm+1u3aBRCkYTaFRC2e7hhJNVFePuLLotfPgr63MNi
t035ZoAPUOtqOHnkkOs/WPE4JbLDJoZaxcsV8bjXTqCX3KnR+7G3fgNcKrzhA0sDHCScqySNJv60
Fil0exom3QWtzeS4t7+G5EZMG47YhfpxIBSqnkJoJbO+iTAVN/YJz65Yoi8L9EoGAhDWglkBUatr
XSk/TbhxfWGclnhpcYiRsL1Va8/OjUgMDYhbTKGusUN+M9uaiorZcNgrudCKuqp8f56QU3kjlm6H
9BBjSq+uNyXa3jcUL5QXiSjaXKBxOKZLi/IeWw3RiaZ7xrwBxfjZwZDW5l8/2vQNetoUb1BWBdyD
XCDBkgV/7SDHkhbZAFawTnYeMV83aKAq9u+gIH30nDi2b6hgOBUtEHVq6YI8TDpNiK/H5C8Qld0I
zZ68dIfi6MeHwAqbKRzRxAQU/yewN1fPARdVtOHcThk+Oq76jxKtUZuqRqAOgWopyHFf/XiLCcJ9
4wv9Oh5v3dt3+UoZnnnYMm1Y84xGwcODbMGRFmFcWXV0X+KfGqAmASuE5XXYDsdVCnwPkdKzgSCf
BM4VSFMHJ/KzWiig1tS/WjeGvEILjLa96wj2xhQaPJ0MRFuXbeXxUFhWAGZOeWADgyqjt4L1GOIC
iw6RH/weL2cGS6kXqAkEN9jnUkYFdDoBYqIeE7TXsqxX0NarloUbOvrg8WLA0gG/TgmNeESmCyHq
PHl54XRHXaOczqWRhVz/u0bHVCiA6oc15lZFb56mKHo/+9sM3KmD4x3DIl1Iy69c3EvIr5inpJk2
aazUr8Ayn+m7Aa1TRR4iuYmotGr9dN6jwwsoTJX68cp9ni0q6PthfrfsJxqNBMRcD3B7jpcl8WI+
+A2Oh9Dmtp4wn4PAlJEFufBEYpbdFxP3u1QV1uNcM/LrZ2FBW8eCDRuEh2TrOqS1t02Afn20pI5k
EneqoxwsuwG2LfDeOyY47bga1Ot0d/LyGwDzlE0V4CJI3ThiqYgLjFOqkEm3Ymofn8EyMKsU3f1Q
yoM9ds2YPdO2976R+9ZSPgfWMguo4hwnQ73XojqP5Cs5kyRYzLWLaeqVZpFl8twarzrixMGSBnYS
nLHtV43B7V3ZqmR3stFjWV2wR/Sk3e+1/qKeah7aIEjXkwfs/NUv12o2UeRSvkce7rU2UDlmtuva
roKNLa/MDgmXLF7T6c1XsBKt39KKcasPhu0d9i3ywRmVZyBZceK2DUhtkJqSZjrYvbyM9WZ7hlvf
y+GjePwoh9NTdKCYFNy793X+4yhMyAVL8GYX+0Gtu5dwOgHHyWYas6rpLyQN0DTHAVQXcnsiPvFh
SCAcoeZEcO+V6C74wGbW/Oi71+2pxuXLlVF+qJMw5cCdoCjSI1N2lw9oIAmgrqbhpGpTz6LMmrqp
ndk9eDZjhfafqBWItWopcsyN4+neAgT0I9eClWJNioaVmN6kwQ7xtYJ8Bufw+4R1PqKHu0vo3CNT
j9MTrDU7+owq2KLZEODD10gAKsXoD2WRny7Gzmq6CxeaAwX8iZ/+Q0oBgbm7VMXEW2d8iG+sDiMH
+cFZDAs8KrBTljRpbZ4P3ukjbboYKmFanPYBxUSq88m+w398ClMSsu4zzdjybYJEaI5cbG4YwwT4
90n2+gSyOsPOdH6je7TXhyhVxe8q46mCoor7yFZ+H807ln9Hlfan2T2uByuP9w4oLZ6dFD8DKMJ/
L/zCLhbuNxbkOR5l0dSJQeAAd4NlYCCV7aSwrLASrCsqM5HshxlYS+7vQSZNtghfJ7pb2Ff8bMoh
gGX79sXhWAbWarox1TvAUgcJvZAhPiqLSVDtdiwuL5R8gOev34PIsGp+ugI5thZxnQeF/5W/Migl
sNjvCB//ndIBz2Vw7Ht2iOApd3U0ARlGsMu/OVdMe1jCkmhPcrH6HwA4DJJJOy9KH0TnhMpFRURI
bmxMqisO1W8vYN6I/VvMfupH0pOMKfw+qZ6S8N2Q30eF1CCTpuF5XnygAg4i4Ax0mVOl3f2QJnU0
IwTWIbgedFERZr+y8/eIzIfpuUH0AwDcdPOxM+GTJPTBQcO7GnCZjqbR71vskK9Jhybq4Gd6Qi7F
/u+BDkGWLyV15OkeOKTcFzzMntmPY3hCcTIudkUNWE3azPgK6hhWihjGchkB/1BtMOg7Qi7o5OGg
bOq8FR/K3OcE140kYYpUBFR1FjhdX//mkQmfrLOSX1MpgBlNmjuv5C6oHUXzLxTqRzCZYxre65iQ
uXEZ+xDkXa0fXuhh9tbGvrc+CZ90KBXnMF9X0Hsma5aAs1c6zodL1heyVziCfR67/8jxtSxHmuza
8bNWF8rYQd+OZyu4PF/L/9cgpO/O4wBoVVeh59QI4O23cF0LpjsCEB6PVBlr5xKZITQR5QrzxPBQ
UuZK/kSA86SNibYht+8QZM9QynkINdH60O/SYl3PAL6Z1VBw4Yl/hHIhI23V7AdNPJmbwUCQNQ6S
PPwbm6HysDCVf9ATLBMPchehNl1paKV7GXyyBcio+5pFmmvuOcwjptcOr0YxN5wBAOMd9Uv10A12
fg398D3N9Wu/lDPxWj3RIlz8sCwl65V6zHyUrPE+9g7SGGF2rLNioqE2Q52ui715OXUIcAwxwcEK
z3opsq4groMzqjXyOHx3JdivDoMCguuUjayc30WRztWyqncRhAm8Dju9Qcth/NacbRWUxftGsKy0
VttbCUPNyHtTpXOlHc4A6loJbQdOw0XKJbQT3sibct1Rijim+AJTY/9NHp+rJ7NjIrQWjzUMuDQi
+HXXaQDU7Amr1QJHsBELo1eDdMrKetvljChJ4aCAnazwHJi75APj9jbFZOSRHQuP19SpOx75aW6h
I8+JBgZZb/6xUzxX8JWfOPwUqJ5GSorCJesbQdKZLqqig7qlFqK1vKjSgYIq6rnvZfAJA4IE6EhX
KI++dpsm/0rLXLABlpXkWEQkLcqx2tzjB41QseIwPkOIUy3Gs8Cr7VxUL8WnWiWW6JbbfsLGTn4x
lamL8AOPxXP/8xcKEdigY8mhRosfRk+zf3rFeebbCVWEFIUanmmEYl45zeIzKzMOrfwhatAkK0+b
JNbkb4eEDYayEygKse6ylzu2554vvWX8YkPXtLV+s9IKGYS69drSu+suP7SeADOSy0OCxtN2nR+o
Vs8stVQMr9GWhQQNbkNXofivouMMd7g2dX3OhvyMBGj+vmescuUQiF76doSpOhOxXIDYLdCy8XdD
03zWrJl8kfqJyky1ts+LwaO3T8l581qz7LvYL0laU4Oe2O1yoZzOjvx9p9LNWWklddr/cfQS4arJ
NXxq8dRfyoDK8UGnDNpII7A0gjDlBoIFu5f31oxjoNc8sYmfPcrcqojhW2BSi0jPork+R37jmX1j
2kqWT06RMWcxEJtMNx/DFLhY+wmkshQDpaEVmRoK9ctYMP6vrUVEiOkgypwCKa/CDTDKlMxFAypO
lnoq2KFFs2PMrJRaeGf3GPi+ko5k08ApYyz2E8pIfnDUW0UtWDJZ80nhEfP+Ukmo7vqM9Y810geA
Gu1Lgata2Ds02EX+kagqX8J6XK6O/IHZCOkbZ95dYC3QJinRm2bSt8fZhWTGse0tVXO0ukJoRJhj
tAwENNeEv4QAi4mlOAlPFftK0waDmMLYVKfv+VdUiRIryksY9/K0JTfcN/jSe+VSYNl2t+CoIc4D
jRPDMAxYrBURQxjsX3BDBm71fRPs4IkXuDXaYL0VLaVrmnGzft4Mz4pp9uUSMhjzRDJ/EsrqQ8Z5
T0hpUnP/ahWSvowbdiVKq+SwXeO7AhZepmRe5hYArAtXn4txQ4QFCqpWkj5lgu7NWW+CMMbANOLO
3YT9djk8YElTiJ5LPm+mfkMjw5nApuzpD5qA16F37kZ3YGtGTLzyKSEn/ZwOwgiUaMBgib3tJ882
1dwhAjbB6qq+rkUfnMeYuaPPfq9aYUHi1+i7imFvihJNzPYzbn8I3RISk+dGupJPf7DFNbjMSdV7
Gtu2Fc8591eDV80pZnmd/hFmBmpD9QJMLlsO6N7XMz9dADTj5S48LIvbUyt/FJ0oljLI3r8CzyQ+
y89SR1irYZKwsfIA+nowJArJS2ChKMMx4hu80a1CAvhCspw9Rf0IkCUNFFAO94Cc+/GNFhza/N8l
xFsZH9YtLyAGAdnbHeqVauMvHEAagx07I631K2b+xc8T6A7v8nywUIpcgH/hjkInYT6FBEJDriki
QEJEi+9qwfp/fJPBDv/RyRsLAuDNm9B6kiXF0ziWy2mEtDtWffC4rd/DVPEF1/5H+4wzLoKSc0uR
Tp3k93+OnmTB8HRdaHN5be8gH6Fe9NPM5U8R4fwK8ltY770iXATDC8fAT8vg0ozZ3pLknfKiT/xt
GG2Oq8j71Vd1XhKScvbLirOZ2ZfcmcWly2scX+cw3uT/RLxSXX2WFGvGfdTxVPTK8NblbXXvwsTJ
8e671NbsQngJ2H+ouUpvZ5NH+6SRI9J1evwNC/FIDn9G77/nrmFilyXq9WFKs418J6xjy+cIOEru
4g9VMHTE2semLp83WpgBRJRsH59D7htbIpsvjJz1RJQm3mRDwh+Rw2XKL1dTrd/pxNyqo1/6wOJS
ZEhyAJR1nbLtYJVghETQBm4/0DwuEFdFWXhyD8aRPIRQKvzOIMRZt0G4nc8rSWceJt/Wz9fGasv9
hVgI1gQSh2aL/VT1W3Au9JNuFmh4doa7orUIja3KGEaOYh92ytZpH7LbVAoZFHvvqGt+B3RRZZzH
m3BfFND2sgmZCCN87VeGvT+4itlskLmhJawEmmE+2FPekBrR7kFQpH3ecH0g9JnzrLQIZN1jJFIO
KtUHYtQieOHACH5Z/NgwH/wgdFrBo+TszXPnCXhWjB7RbHT1AEIeYkp4HZ6/P6Xya0kpV+JYmmYo
shxWGVITEKSfBhqEPXxczpOxN4j584tSiCec2R4XR+EMYgxJPY1LS7CbL2dZf5iqHg9hBGhN7LMY
2F3OM+pM28DR/K7RerP7I5NFzTBQyZEQd3B/rcHwFfzSWVFVfVeb7UJ7WTEnH0bS9R7ggSpLMTfo
ZCu+TqTovfAMBWW4uiYs7IYRfMa3QWWu9pf45LWzYChTTFkpbWIO2zp0YRGJZOvaxJXkf+lffJ6b
htE9O6yFKpLwFP5t2bot9qGESIqE52sgouSDZ90V5+6c+zPLj/W8lgpepq4zJbfqR6wbK6Klg5oL
0LFiCC89ghXu5hBThvCpIKt1s75MxYEi/GQVzJhqo3VVvn8ZJC+TAjY5kW+0O2/xXWum6kb0rCVr
JmgfeYYPlFMDu/7M524gdr81N+WrajEA6zbvzd3MuSssfE6O7WhiM/bTlGWXkbUebtgRapdhrrIb
LzUhbnmZP5fXMAelVchnHUyl+EUQe/83m5Ara16u+mQtktlITR9Es5xzgFAv/JCM6GF3ccpTGIT4
ZAjvFVye7vFYJ3RgA0QR+2DXm/4mj3g6+DvxKKlNUbwMEiAtgGQae5VyokLcdtTWA1i20r/5+LRM
z0aYK5xpjdScLEBrs6XPGsFhipK/nuul3nQJ/vX8GokRDgCZFATz2yJ0wH1PRxVl77fgnZ+yTNOY
MMxArfviZgZBxQgP9dNZKvIyG6T1ZwHayP20GqS4rBuIjbGob/0jr3CEI5+n3OYO1k9EKl+Rawoa
z9fPzY+2cxi6Kp5Fan4UPp+GLf2vHM95nD04yvnsuwedUCYwQuQOiVcXnO3xWDLmQnlXNdenNirG
+ylxJxuMZh6jL3QZe9zNS04iVDvKtLmmJ0y6fTvr3fEkvqeeR2lWYgkhqP2QK44vkp6Lwx4fSld0
PLKDKKemPF2zBYadh+QJnl9YNQkCi63S8oZCNaYqgbHdWYypr3Mv8y8gXkIjeUtncKaTd0NS9AXe
3ygqIYe9QMu3K43MVANEiojXCpkf8tIvxMbxKqGHjYkD8MDTYMd2QhfAiU3zRbnvFegLEg+CBwHE
OPhOB3XWJ8wm9yOVh9L6tGkvwBMbVW51qDXjRYL7ipsWV+bvWzpDCWpIY1Pf9fT6BXXNyaWq/MUN
AZ3sSFWl8d1tQP78MJ9q6znUPxxsQkYI8IN3SnH/mbhs2JuzouBvjS5attSaLkOkFQzM3zlTe7DF
Kea/tT+mmHTrJKnctuE3Qi7venHseXhYFQsUyp8c3bjzPKWxwMpm
`protect end_protected
