��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���l��o[��ɴ����>�$��	6������b@�	������b��VJ�o.y����L4���Z��1룠������	�<�~���E`��-�R`��k��-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_d
�t!���N�S��گ/�TNM{�C�5���M��;����L�S�:�{���\p<��)�0W��B�R<Qt��Ԁj,3Ӂ�v��`s�HW��眣�U�Z.͓k����W�z�N��VXi^�p�ޒ�}���C�U+F(��o8m�2�0 ��r)Mo� �R~����u����}F$�|�,s4|̍���W>���%��wE���*��K;�p�����I������R����{R�����n��A��[�͛Ϻ��U)OR!�<�O��>W��j�l�-D��D;���j�+bq5#�[`$5z>6��L��W�C,Вy�4n{"p<��+��JL����g�'g���Z$��a͟�@2�H�wj}� nDV!���B!] �8+UsC��癃�rM���>��5�ƈMe��H뛖�qA��;O_����G�< ,�XL�v|m+Sg_����?�)nOK�78�l��\ad6C���L��t�Ĝ�u�H����/��FWx���m�c�gR��|l����C����e�	3l4�MI�BK,l����W��.���zE����U��
�}*��P�]����<_pB�
�ϝm#���QD޶��E�����7ha$���s��J�3	]w���8M6�I���� -� m�F��z<�t8/z��/z$ɉ����M�Fa�>�]P&���&v�P�Eτ�'帐^�I٨�������0D}=�Q����;M�,�푄<������$�q??� 1���߂x�$�Gk��@�����v�����_E���W}6��=eZ߰b3͵&�	E�e%�?���A��< ���h!�U���$���&m��Rti-�Έ���$�u�,tT��
���t�����q��l��@:��b��?�N��w'�O�0���
���oҕ5c��l���/�x5�鞱-I��>Uϭ.���[���7[l~P�k��i�`AZ��)I����^Џ�t)�rom��!��>�sQ%2%�Sj�c�b���u�Y�P�,7ӑr�(�ۀX�/���r����m����LF�_�t|T<!��G�<qis�*�gpk4�jl�q mԘ��p����������N��[��i�y����X5��K�+�o�ZxL�c�F.�YxXu��Nġ;2|��G�6� u2/*����4!l堮9��8���2h
�L���1�Nc�v?L�<	y���3yT	��D����h�<w]��Jӝ�AI���i�ᯭ��(s#Q����@N�N����"wzp5]K��R�G
��!�Si룘g�MM1%\Z�L���0�c8��bG	vH/t7�h��.'���yڳ�@ԪخIќ�)���(�t�_o�.�挒rӑý*�RnI��.�㨮�[Eg��Q�EO��]��g�4)�Η.L48ђ��}Tŭ�;U��z����rk���6B>�+Ͼ��YEA����/�|����Ӿ��r��N��1�����c)%}�tr8�qtŘ�()ͣ�`�Y�O&�V]����1k��ό6"��7���ef�G(ib��e�a�c�|��E4 ��z�XLF�	�X�ss�R(Z�.~X�H�5@�������7��7j/j*%]ܴ�ާ�5�#����P�ÌU�1�ʔ�.�Bљ�ٛW�$�W�(�"��nK�oV����/�������/��*Ղ�us��Z��s~m��B �{-,(�H�Nd55�C�-�g���y�Y��1�a���������(e"�"�ɖ�|H��T�a�͛��=���b�?K�u�>�,F�!���@���|�����V�1����<0�z@U��ML����[$)��q�H�&�=�6��D�Q�� 悾�QŶ�C3⨒�`�Eg�Ҡ���X�K~����w�����''$�~����n���}�!�/�����o<��޺O��1_�Vڰ��e7��t�'��C�p��fPc��J�� �Ւ��ﺢ�n�L~�6�ߒ���������:A�/�w�F�Q֋&U���)K+/`8�?Wbb�{T��,�GhZ�������?��7ϖ�V��׸���Yծ���L�B���)���2+�/V����>#�f%Y����ɞPp.[�3J'-�%�,4�?�����r9��˘ �MxȖ���2
�XAL�]�}��,��l�Wa	Vg�º�|��f��p�GB����Q��k�=K���X!)&��W�HE�1�m�X�<��X��3�Z�=�,��K�UպϬUf��L��Q������}�*�k��36j�W��L�"6Ɣq��]��P\F�5J�$6��/���_M�n�̻��i�O��,O�Q%C	ߙ�����U�<U2/Zj�c ����x��k����0$�o�l?���AU���3YŽ
�Δ dSgc�*����S ��,��9O��w�����iS����.=08&�قB���H)�x�_0�Y���)�>{����2��x꛰�Y�:)!���?�M�U!�}��������ؽ�.)����MK-��>?R���H�s=2}H��Z�f�!���G�R�ս�}r���]id�
�W�QS���tV��y�E�׋�
v�m��b��]��P��x��)���j����k� ��7w�5��k�$��� �P��Z�\�X��d���=���)O�T�W0��R��Ё�}zE̜Q�՜,��2\eW��Kt��u��Z�k#�%�1ڐ�_��bDN�t�Y1�K�񾂌���>^
�-�Z�~�X�4+�k�i��S�{aW��a�Z��E�Fπ�:�"&�ѺN �L6��Ŗ���q�SϹ`�V8�Hz��X ��р!c��ߨl��X�_2&*�o ��p��`\	"]N��LE��m�H�J�&;W�t�J|��q��E�e�Gʪ��ȫ'�d~���E��]KR�q�!h���W�	��t�A��	H�:~'�FV!�Gte ܦë�2��#�7�~�Zp���V��*^ʝ�/<S��|]ˣ���%+$b�>�U'�ե1���u�%W�]�Z�Bg��9ł0���^���fZp���$1�X1mc��G��jd4 ��?�L����	��2�M��l�4l['�z�P����a�B�2Q��a��6E����b�L��9������!KP��J�"�Q���jm�?̺N�c��7���g����mދ݈u!BoT�&�fO�V0\�cva�S3¦��y���锽ʬ%���C)M%� ��)��¤Ss9%M�}f��lo�oo���������+=���t��iyٔ"C�U�
Yh�)>��4��q��r8�jrp10�Q����:�-aɺ)���)9M?�̆N��,m���o�z@���'q�I�)���8n���Da��F�L�Z<As���a�52��bP�S��:dR�V�k����]�5>ւ�+�]�W�vΠ躏J\�R+�Cg�:Kn�����A<HH����)e�]��g�u��L�&�a�>g��R���)	>UgI�k�W����#�h����jjh��nٰ!�jӃo#��G���~��S#fhH���b"�u7̍6�p�* zEy��9�j$�͍'u�
H�t���	���e�D*`�P�����T�)5<��ф�E��H��l>K���b�|�У�����K�f����*�<��I�*�WA�`�3��t� ➄�Z���3�Hy
��I y ow+-�+nI/;�A�,*�z�maI;\?�$/m�u+,�3L+$J�I���*>]��B6����.���[��
����}��㥩+�vF��|3 ����G�E�(R����͕0�U�E�fX���AvT��1�1��I��#��xg0{�NUx���u����p�L$���G�]E�ip��-���|7g��,ू����ɧ�a�nx�V?���f!� ��\g��%c��?�!�A��A*|�r�R5>(>�/��:K�1_��	̪��l��?�h�֪|)�����Ƴ7�6��%ky�p����39�D�%����R��~����`��@�'`� ����Mp2���K������v���2�r�-pY\�e����m*T>o��5LzZ�[�j��P���ˡ8bZ�q�{۬��L
�B+A�	"�9V��cu�RU
�٣�oh{O=8��T�n�S?FQJa]��CcrǴLƃ�����.p��$KτL��GR*瓍%;g�6b�v��!��*��Z)tiy^���'*-zNB��QmC��|F�H4��&�{yUy�2e9�sk@X"i��T盗��Go����?���1��@��ˠ�qt��0���t�l\*7.����ȝR�l;A�՗���]�]�%%�@<$t��E�zy�9�;��}{⟱��v&�"�X���j&��jT���M�	� <�7*~�'XK���:T=��a��# w��m�<��@��"�g��TDz�ֈ_�X���g���W��ފx<%��V�r٬���N���S;�𬔆��u��u�ӈ�!�oXy��M�槻qS�yG�D��7��~6�sM)�����E��դT�F�#pZv���hG<r{s��[0�t�)��X�<RJtN� �5V����e���.s���ѝC�����r};��Q��rw��e�忝Zb��DS�q��+�
��A3	7c���ϩ�j��F`��U�X
�58UXsm��ֱ����uL�)�C��ۅ��ƠB44�|�7�A^����T1��P�{$a�JD�꿧�����FPZ~�r��g����N9�0w!��� �^=^������ԓ�N�����>l}�n�<u{��l��Y7I ��y�0ޅ|�O7-��W���B�|�)HeuM��<�\�!4^�����rB#U�a�0��g����ܐM��s��K�c����n� ������{t��M�3?nJ�	�ˮ�F��w3�x���u���?���hŎy#HLrW�	��q�4m^�в������ig�N5(9�W��ќ(�c��z������W�i4�(��
�MU���a]ٶ��T[@���$�@��V2݅��g�1܃Դ���C�U���DZ����u��c�߹��r���{��9J胷�I������ �(P'�&����5��Յt1`ɇ��z�V��DQ��
��j;'��s�wWB�UW��W�y��?����zEЃq�K�n���������#�<���pp9��[��O*pq=���eL���K��Z�϶
̙�-+S�Z��t+?�KW�L�K�BL�DY"�k�����W�P���-��D�hI.z@�/���D��޲�X���H1r��w>/`��2M��8d��֬�����ŷx�'�&�#Hc/�q�]1fm��pQ���p�ש�l)igY[��Ǚ8B,�Sdo>��'��g����w��Z�;�/%�'�=�Uv�� 9D�]Ym��[�|�x��4�+'Jqwk�i605��B8��S�����A���:�y�Ҁr���3�q��/I��Jg���:\p�K� �9�8Ε�'������s=�RATVG\�� ŏ�?�P-|��gޅiG�x�}Ɣ4��"��t��=X�e�#)�dg{3��=lfQ�݇����/��EfH ћ��1����މW�Kj:�d��Jڈ���u�FԌڸ���#�q6��3���Oﯫ��P�ǥ��"�����$���@^���Μ�oG���S��B�HF}����=����*S;�(��֪#9��[צ�C$�s��qaW#�Jݚڬ��7o��E"Gr���k�&�]�� �(�.��ۧ�oQ�7�l	j���AV�O��|�%$���^7F��"7ҟ�S��
B�N��Q�~��� �'ڼr���_����c��ڧD�,8Ő����RH���T�8��I���N� W!�jo���zlr��&�����(u��e�CG­�ٰ.3'��@-�;�Ȓ�����^V.��/�����0��o��9}Do�X �����f���ٔIj���3����u�Ap�)%��8~��s�&g�����\��s���J������b-�z�Y1�Dx�S:�K,I^9h���p3k�^ˀ�ԁڞ����&@vU>��[�Z�����{�1�;���Z�� 2��~���D`�`�AM�?����(WD���._�'�3,@pS������,r4�Z�~��L����mbCh���f:( 
8���A�T���g`�2�ܡ�����<�n��#}�Z��A���G�c�S��W��E��K{�!Yui0�6�&�̅@<ꆐP�"��|{��G��ql�ucT*2�=3�7�"����YQ���G��S���������$�RӲ��ٺ�����$�}c�Zo����ol�x�¹A��R�����:�62Μ$Ye����WRc���9���|�V1�P�ٓ��l][>_S��x]�7����^�θk�P!�ZWA@�f1k��	���6�/�K��H1v��H�&�p)YY���|b�Jq���S��]K���7=�$�Ab�l^G�L�Z1h�chP^�d Z8��D�S��m�&!V�RY�V��a�S�_�$�Ї��aЧ�L��oF��Њ�]5���*5qB���N�4��{��%�o���G$�n�R�`��'�̉iA1���WI�8���g�A�$���8*|����%�����%��M#R�+G �V�Mh-���p�԰�>�i��Ətϣ>�����G��~���&��	$�&@�Fǝ��?�����A�y��Q�0��|7/��	8�G^�e3�M��O-�d����N�rw�)8	��P'��S�ͫ������a6[�����RE�Ҭ�  rɳ�|x؈��z/;�~�=l6���{��ǯ˙�a�W<�J�L\<���?5x�NgDj��'�wO�vЗp�p#:i��[keU�{�,"���Ӂ�O�i�`��C��vf+��#�^�q_�LN��>�J���U��7{�;����i���^�:�$�1.G���f�8Rjtb�ל��@I��	3)J��1Gd�n[w��*>�u`Ro��ݔ�n�������j=������a �pn��<�=��b=��!���w��O���s�\���?�|��ϣ����Z��g�E��x#g4�uw���$a���H�b���X8v���jT���KU���2bU�HA�+�v�':��q��4��R�����لbD�t��8U9d��E��\���YqF%��u8�U�%�Pr�x�\b���-Ek�J��+��nZTw���l��3lJ����-GO��p�*ά�7WIˏU٠�=K������$�'�� V��c�MOP�s��Б�i*�au�k��T8��V"S���=� FM{�@����ʑU�am_�6�+��%��3��Z���k��d�o��u���*�N�9���Օ�w��?
yp;���re{XO�)�?�IϠذ�.��:* �(C�	�'��c~O�y�%��-Z�6y��ʚE�7�����.W��<�Ad� ;�����oN�?������RCk��������}׋ZG�2uS�i��4:*�d^�6��G#Ƃ_��V#������N�0���5-nm��4!U��욨g�y
��0$�>P.�Ǻ��VezE�#�W[�}��/0���>}rW���lZw$��i"��g�`[xj*f;�Ǆ�e�'�����۷E b��Q[�}�,	YY1�Y*�(#�o�aKď^B"�ZiʏG�����-�4�!���S�d����Ap����UF���Xc�5�A�~��y.��q6qK�-��$����<.'0]��Jq	�K��*+�V���bY��,�����(t�e,��E]����nRa �a!�紾�n�{x���%	8�����'�'� x��6*tQ����-X��h,�jβ���4ݹ?���f�Pc`2��<>8r����".&[rx�'�L� ���Ԗl@�%������wý�{��ٞ-����H��Eeΐ����>[�(��*�79{�c\��ِ��1�+�����PZ���V#X��-�y�`��0
#���/	�<�^�*LQ-P�6�&��_�==<\��Z��>�*��35P��'ZGZjѩ<VAoT���5�"�)~�N���x9b(mV�yX#���F�����'��l��
�z��8;/L�^F��p�>1;O_i����\	���ж5�c��ݪ�����ב �D�p�p��1���BU%�ط]eW'v�^�LE�d$9.�f����6�L�V��0v��$W�"��R����:׆u'a[���vt)ku�K=�7�w\
��%���E�آʠr��j�a{�"�/S�,������*�o&���g���F��%A�w���N��&�NAe�H4?uZ#f���H@�a�tΧ\%Qny	��`G�O��'�n�\�S��o�NQ�t[r^~y��%���kO�5/>�	�ZY6d�Sk�P0��:�K� hGl�ȼ-^�zDi�����z�k&���K��X
���T��:��@����Eak����-�Rtl#=R�
@	}bg����;K,�c9�}�#�I@���Q�W�`c��ScN�p�l8v����{]V}Դ�.�"Ed].��u��;���m]��2���~���,�����hz�)#����@����k��#4�\��f~��p�f��Un9Zk�J5GE~�?���{DU��]b���	�T��r�Oeʠ�劉�?�h|$����`�09����)���*_�'��ݨa�K��?8H2T��4��O"���e���0e2����uV�6�����0Ÿ�jv��^�r�����}�p���:m��
�������U�%����uԲ�k�C����ۊ=���J�zY��Rf
�y֏<����H���O�����ϕ��IYj;9j�T��כ�z��ZR�6�`�E�4��}P0n���%��
�D=��g�P��#��;I6��?�hR��,�:�=[��<*j������H/�=�$���{�z�<T�h�������v��R}�4��mj`U`(�ZX��ZC��G�z]���/5zB�>I3mɬ7j�s������<�!�a�}}��� �D��Q\�:%��\���x��s�P�	�/�6)����5�~��u�� !����!��ݲRܪ?��L�g��1ڂ_<ӳ��,|��~�V-��O#��+l�Q|�m��8hsL���೶L��x���`k֥_�H��)
�R5�E�ӆձ�����>�()�I)oSVa ~�OLi��3E��fCS_��#z&���ɤ��fE��D�6�xc�3>Vzpcz��M4�`�5x�rB��ԅ�%64�K�hN�)��s8[�	A��jf����n9f/"�J_���ڤ�����������9z�_����^%��Oq(�v���O��]��Mڷ>��"��*�I9�u�&�8uv�{�%�����8�k�#�p�~~���d�ȼ��Z���t�o���4���F2� ñ�:G,E/�ݜ���լ2�	��D��1��g�~g?��`>D����}P�[]DR!V�ҙ�6�������̪��P��;K�-vp*�0�f캕W��Đ0�|�'L8vՃ �d��Èkݒ�ޠ�]9j�Ǣ�d��:�}]ˣD�n�֨MG���۳P��X�vUť��:�RJ�!:��m�?[�d-��rf�'[�$�ݪ�.N�'��	οH,���oV�4r%��ޏ��Z�/��&/�m��Lz�`E���X��1NK������	=p'q��xP:a����/�y�י��<"�s�WV!�v���J ������/jU5��z���.7�����\=mL4̢u��:K>ɐ:K�l�q�_�vo)^��V�2���?q(��m7F�~4�Π=��ە����I���CZ+`���haD��LI�ա��T����'G�e�eO�w9!a�ى�$ͥ1�wf�D��y����D܏t����'*K��	Sw���:K�M��t �i�5TܦO76�����s��9}r�rvM�#�q�8z�+�]�&�����C��ij>e�w�1B������xȪ�E�Z�	蹇��_������dKs�V�<=���q~�F�/�]0p
�U;�c�BY~��8�_$�0ff8|�b�6p���tB���%���o�w��m6Xq߶����9]���ǩ��V��&s���Sؗړ�+,5׊p6��!�w5�[3���_�tB���RYU��b�8�&3=
9��q
/nK�CW�#��ҫ�4´�)�X
N�tD4[��<��л���M��Jr�$��|I7�f�QwKw�M�s�������֣`��]��UK
�k*	h����w�%�o�=e�|;T	 v���������ݻ���<�!9��A\Mq�-�)0�����¶�t�}�A���������ű~���! ��ж<% ��7IeZ@�aE+��]���L�Ό�^�2�[�žA�u�
�"`�3	V��{J� ��Jb���1|nn�9�\������9�r�l$ɂ��&]����[
O�妏�WzR*&��-�s�P'f���b��K��.B�F�)\����}pAPhc���`jR�,̫|�q�-/}ryߥ��Ѧ�F�3yn���CN�9ι+ �1$�aފ>����������>��T9J�-o�Ǭ���A���?�E�5=���nb��j}u��Hr)C���.� �^m�\&:��F��m,w���B>T
���ŃXG?E�������є�j�u�zb��*�eR���2���٤��2U''Wbl;�3�6{ű�AbA����qp���GD�wJH_C��Ι�'��	)�5!Z� 2�شLl����%�����_)�Ն�C�3�j���:�%|�xr��X�� S
i�#���V��hj>T	l����pΆ�	��9���x���z~h>��y���
2����9��o����A�Uw�ugCd͋�X�&Q5��|X�\
U���" �u��h��-3�ڎ��/�2����H���e(��t�}��S �+Y�9L��w������5O@�_������� c��./5Sv��]:J>zrF�?E��i����,J�k
�D���6g?�<3��Ҳ��`?h�2}��yg�}���.Aw�;��Pw��f�ǆ
k��*T�7dQ�9�ȇ��W�(AH�y�|����C��@J���F����Gކ��㕞��nL�W�8��^Bzج(�J�D�$�X�,�Ŭ����y���J<�:��5�0�y�B�}���{���l��C�[�_*��{7���U��`{9�(j�<쯡�q'^�9���*�Q/�s���Ag�J�駤ܻ���l���ń�(��7�wd*��A	��.��qf�����b.�¦m����~��<88
�:�W�|M�NE�D�,[���^�]Զ�k{����!�S�����(���{�ok@�E�ط>�0������ӾF�r���f��gNP\��ۃII!u�Lk@�5
T�r� Ⱦ�L�X����<ߧ�3^LO��Ӂ��z�k����.z�����S���۪E������y�b�hK�ڂ���w+��ǌ�� ����̋H3D�������^�M΍�3��	�Z6�1�j�@&C����\��HL��V(a͑�����w>'���P��*E7��֨dHa-�O��O�pNO_F#�,��+Uܩ~z�ⳣ�h!�
so
��V]&tõ5T��vM_g�&�[}�iנ45���!�U�,m�T�z�N+�LVJ _`��a&
%B��Y��	�Թ�H�s�A�nT����2K��q��L�m�'	�Q�l��Xn�d�WB拝�:Sɭ��c��v�4� �����g2�c��IR�Ea_l��5���ȖVS�x�~qæP����r[�0��P�h,y[83 ռ�1$e����e�D����!b2r^կO����)��ʀr���~�,~��E��ro�-=@V���P�e:P�U��)�, 2	e;Ӡ՗ki�j}P=�k�:Y6V� T���V>�C�#d��ZJp�s �5ⱍF�EQ�!����2�\��	�� 0��X濧~����Xy�-���D��V����_9ݵ�1��f	`�Sv��1��j��B��/�d�^]B��p&M[����"�n&Qj-@��1��]|����_���Ms����Px��e�f4�e�5����D��O� t��9�)L`�S0���O���@[�h�c9�{eqPq��#���.������V&e�~a���88$�Q�����w�_B�v�����S�ˠ�V}l.G9���5s��w����N�y��-�=$f��w�43��b��+T��=y p/F��JI�:������X���F��set�p)�ֹ����>[���|���*�â��~��h;k�-:�j)��������shi�ŕ��þ&�h�P^zNg!?�&�,14��]�6ڿ.+O7L (U7�vf����C4���P���q�Q�h��Q6BI�?RW�_�>=�XO?��;���� �QuR@�1�ټ��5�ge�^o�z�$u R(muE�f�;ܾ�5���� J��d�׶�柿q�}:;&5�F/�T�-����Mؠ������g�Λ;<����BI~Bj#���9Ʈۣ����0��Xx�G�c���O���+m�D���C	���Cw@ݩʱC���9�N#@�Ҁ�In�?Ğ�U�,��ʧ ����Vi)Vd�}�<�Г����L	���.��9�@0o�@ k�$���sX��X輭d谥˕tG��	��E��)w9�sue1��y�"QN�
�c��Xwv���R����UJٳ&c���(�$@pfj��4~�ةb\������z���4�Ji�%�i�ʸ�H�k�X������.+,����q?�,��k�Ce�j[�*�E!�ZهtP'<á��af��Y/�ҹ�[]M���8��hE0�p�'-�m���܂`֢�#5l��|q�H|�f,�V�-q������,��5���ݸ�BqRmV�L��`�,�H�t�����L�V}⠳��M�/��w�5UG�?�����_8�"REq��Z��_y�{�Ƭ��}ݸ�us�0��B����K�����>���D���A9��q�%�d�{��*s�-�*���j�+IDCG��8[���a�]Z�� }*R�[�T@5z&]��
��ΔZ�4*�6�� A����Lf�
A�@9H��d`�q/]���_��PK�6��4��y�!�( ��}0�^�O���N4�������K[$���A��-&��%a�3��~-?��$�f䆤�)C��͑ޒә"pm��/yb�4P'gn�Ly(|�|��,��c-�sʞ��0�\�w8��9Z�J���y�,z����|��:�'�0!{XL�_�3Q�l�{�+��S�ī5�����O+��]��`+���C1޳@��.�� ����X����QC���I�=�V	b27��G�Px�9�?D��Q��H�/���3�����>0��-���=kx�N�B��.��B��.�~��p����g�+��9�$ n�)�f��5�.Rr��M��	!zt��MS� ,e�����3�I%���i�v,*�9���77"l�e���&'�.J�h��!�B(Yږa����	�/ϥOf��%O��͏�$��*�z2�ƽ2yd��q{���Lu����c��n��<�8ts Q �!~�lNT�((�`��15:����L��鴺�p���q�\�U�0�1����wC�`0����pݸa���iO,l�6Q��*�~�TU���M`�!6�W�9�H�ǈ�v��I����vuN��bq�.$�jxv��[0$cx�jU�0<zp	_�5s����)��X߈��Db	��)ih&�[��G�f8��9�k�n��j��loyXt�170�L/Y�"�]����?�1���	iF�{����-��m>c�:�]QKf�z��5%��梪�.���^T�yAiof���Az,&��'����q�օ�Fb�4��W��x��¤~�Qs/�B1(t�<�YE~�$�tG�vݴ���������'?�%@D�,u����p84:��ݐ��5E�X*�L�W1�G@�L���(��"�M�bY1V9y�T�@�<����ׅ�s�B����"e8�X�SP��,� %D�yӯ�EOI��rӷ�bs�[I�0}H����s�DH�y�x��կ�j�w��m4����ݏD��5�8���˞����@n;�<�Y��d+����^�e�P����B�H�J>�e�p�q�����h�L�|��8�X?*)����!����ƥ#s�95#
��˰�d`�1�͡bH9K����`)s"�/�RC��C{���Mt��|�������D��И�R2d�g��9Hqp������_#-�9��Y��$)x��5bbC�m�4�'��4�Uv�68���.U�5��ؐ%5�))������8��F������*Z�4�<�!l���T2f �� �D��o��¹��9'��$��w���@��)�C$������'��q_�IO�9��Z.�v�d�G��>�qS��Â������������o>}���;�*�e'�'슿�7�1~���M�X'���uZtuԌ�x=�-"�L�(��V]`���z��-�~��{��[W���|7��^Dg�?�r (�?39G�\O裩��ލ��C�E]�%r����!���xƴ�!�����{�1qn��Ʉ� �{�t�(e|Y���h+�0��J��8IO�9��5��� û
�;��A 5T��C���Yp��H ��*Ξ��)��pb눻�$���7�R�ڀ�i�6fI�7}��/N���i�K7�-�HH�5�4�;������x�<�hI��Uj�t�WI\Xs��h~�����I�faR���;���(Z���e�!F\����[�ऴ��3�{d��jB&�8צ9'~�����2]3�b�"��3�0���w	M\��YlvHV���\�� �BJ��7`�Ϙ���Cs�Aq�-V�לG������' �@��	[�-ͣ�l�!��1��Q���_��C��4Ȱ+V�����-{Ґ��AcN~|�ɎP�hFL�ë�ڇ|�J?�:��t1a��}�	�c�CJ��m�_�m�h����ǣ��:P��E�"�ì��\D��9��E���'̑�	C���q�zZ�^� �T��i���iv��<T5��C.7ϔ֣|��G������=���)�(�Wc�v��]��C���p�D�D�=��U��|Ϧ	B�? ���c�m�B�̽�0��y|_���1�^�F�*��FbK����1�������Q���~OƹϬX.(a{P�*��Q._X�/�ɦM�W1�t"Ўo���)\�w	�qª��:o
��ED��%�l��qE�B���p���W>F�{�����8���^o絊A���>����}�}���H�ys%��5U���	n�e����$&7Zǖ��s��ܻz�!�۳@�:��#7�-����1_�ST�
��t"�ׁ[�%[!m���y���;ܙyt�y���MV%~Ju���d��l"�Z���#��٘�o�V�
��fkT\��
0|n�"�L���j����y�r������i�v���E��y�%�2�Z㭂� �fp�����l�mF����q_l�p?�ne�ɖxRW{�&�F��g��K,��a}!/|�&q�\t|��<[�ٹ�Ġ2����Ս򬺀X��3��6��j�H3���M���4���7*��zr��8 ;T+-�T�F�(>�^�>��`��G�ovEv��~2@� M{�(�
��7���画qYJ<DX+�0�,e�".n�Z @Ҷ�Ə��"�t7��A$�E'j���7�w�0��=��z�[k�]���Q�~�b�?��T�#��P�t���g���iѷ7���h
/^<���HU�\��C��4v�{/0�+1��=K7�}�[� �!���f�Y2���DU�9�Vs��&%���V�щ�X$%�yHp���Q[7$;���\��R�A7��2Bw�z?>\	0�&�/�����`��z�����q���fͧELb���;\�<2��j�)� �Ӿ8�0���ũ�������!���#�~�f�c�Z>�D�� �<�-y�?�I��˔�$�~@BŽm5�|7ȷ�I�^˸	Hr����8��3xޥV�Ҽ����C���}E���������R����V�=Gg���׆�ڸ�8�h��k�Hf��:AN���h�s�-�8���۠�.?`raCբ�iY����g֨�mHu�9HS�T�ha���AH��e}�#h�L	��vU)�����{{W�h����eze�b70���z���%Rs����pW%=>Iv��P��a�IR���b��o5�f�N��nR;!I3}�moj��:�c-����)��~�jki�$���`܃�p�٩�M�xM�����4��B}��1)B��n�����"����?�Ǆ=*_��,��X|U��AiR�8N=��&E�O  ��ʣ���͕.�x�� ��ID$����~�n���%���msN�)n�R�.�c��!FO�?:į�C��W� R�:�= $�l�t�#����z�<m!?M:W�#���t�x֊� �r�c�e���	"�������] ����%2/�z�N'�5>H���F}�~��E�ز{�NO��h]��*�M��c2�sP�y!�5`� e^=�İ�����$��t�r�ƅ��t���nn/��;'	�f�^z�����T����C����ю�lK��v����C�u�6|��B�?s��Hoa����g�掑`�rڳ��b�~dx��}�i�Ø5��iE; ��D�z���� Nv=`�������?��
.���c�֔L~iBÛ����	3s�n���R���A���S@ ����D@e�(X���C,g�7��֍E�`Qp1��)��a�Ab\E�{Ǎ�a�#2P�'9^a�A��>�XG�J�VP��U�9�j�Wur���ۯh�4��O�2﯁��[�+�}��Ўf"�ݸ��7�B N
�Ϩ��oC��'�p�x{];z����>Tq�z��Oc商�/{X6��p�����#G�$i�lD�R���7�+��S୍h|F#�M
з�N�,�SJ_o�{�
�Ϥ�!ݭ��2Hl4�y��?# �pV�ݳ����z�K.�Ju���rl����ɠ�|H�q�M�y ��)���o	o�yֲI&DI�������MPM���lG�Ku)�r��͏�1t�7�RI&���/5֭��ܢk6�M� d�Ĥ0V�������I�T��I~��?�Zk���­x�M��ABM�(�\��u�*u�)�4O��	���c�1~q�Uc�1:$�6OWG��:S��ǃgd-g�w:�􏞴���[�SK���=�)�pД6س�̳�q����1����g�V��Q��J�(��ZP#H�B�d*HJs���&���b��+@����� ����}p��U����r[@�� �����ma�������=��B*t�}�rV��k��[�?��:�B�g�I�(��A��YjW���@�Yt���Cd�� z�Ꞃ�>R)U�-r�@'l;����pZ��	�Rz́��/H��0`�~9h˔f��:��đ�O2�6!�o�"�����~E�w\�ּ���x��Ma5¥M2�KuK�V�� f9e;��8΀>D_'� X��RȌ�	�"0��i��3���h�w��E�民�8
3%�1�a���U�y��.�>�C�'nk�܇��/�B��J ����k|�)p�q�r���3���tԁ�ڒ�(��<�;�����G&.DB(�y�"?�F����2߽��axJ��<�CT�uY�}��N����K��?�{l�C2:��!8���I�8��g7s�|A��-���s\#���a�Z�A�uBcَ���:����*_���Z/T�P^~)9d�#NZφ�I-���V�Ӓ/��U ��֡*(������
���Ly~��۷�z�b�!D�*r:��Hvՙ��$O��]5��k�W�pB�0��d����qT}k��&MI�7QขdZ�_�z���ew$y��.�|��ά!���bϬ��y���N� 
���Iν5���Ŕ瑓�B�a~�3���V&<���]On�ې0Gun���!�%�-���6�p`��j�#������a��@��}DHW.���J1y1_�Z&Ng�W�Gdqg:=��Ba`��D���.��J�⚲�Ri��IE��x�|�u�V}�p�Dz�N�l�ǧQP}v��e9����2��h.�N�D���ܲQFnP-���j0ַ���h��T�ྕ��+�IN$�4!9��I��<��$
"�ǉ�*�9C�B1��S���ri4��=z�Ì�܈��e�a��nB�Ln2���=�!k����7t�h�eR�ޠ>��BfC����P�W��K&6�3���g�2[�+�LD~f2</6i���ɸ�x�F�FyΔ��Z��K ��q�d|��PpԆ�^	�����d�5����k�d�H2�B�'�Y/ ���������dX�qKi���e>�������w�m��>���\�%��������3k�!_� J�M�N���%f";ZSV*k��#ɋ`h��-ܘ��½.���^o�|[������J��X��%�\!�%����Zh[u�6��!��.78��0*7{x�C��)�׍�_�yC���K�4��'Od\��SxW��`R�	n)j�r�9Ksp�����*S�+zb;�׳���,q���:Aa �����B�a��0���,4�KHa��mG�f��uf�*��k�lVrQ�f׈Jz�/����ck��h�u��������f�tC���-�;�=҅���6kȅ�8�4�������oW�x��y��\Z͚}��d}�=��\0���k
E�}��~��&DS��d'�o��0 aR�]��R��8����Mu~=Q��}"��1�u���l��z�%dBϛWR2J$"�(���S��c#u�W�����(ӊ�m!�t�J��]� ��m�� ���Pd��2��'�ʵ�L�!���Qj�Z����' wZ*b�B��ǣ��Vv��3|p��O��,�-%�`�d
����q��J&S�mҏ|���uu <.%S�3'+���O�����J�������yx���������Z�a��CfX�`�9��@
���:�#�QZ-�Q���t�'�U�O�����끷���*t+d/�#]�K~��]�\@ֽ��ۉ-(�?��Uc�A�^�F�f(&�ӷ��ͦ(���(y��+��X5�k�ߣ���e2L��.1��� ��Ҡ��m?�P�e�p�<!�o�nRM�1�����?���+}F�a.��&��@]�FA���F:����6Bw<L���b5���@(wd��b
�ɺ�A�K0xEJ�k	�\�F���&���J(spN�zxk>������M
]:������%�����--	N�z�.��4�T$���ᒽQu�H@����	�8����!��������FB֨Nla���<����6��U};5���������B"�g�"�Ha܍Y�dBI��H�e���	t���0�%�9��y4�l��� +��&lu<��~b�-ȹ����+P|�j�%�R��4�i��\��V��nm�V����8�K�f��0���8ձ2����FU�Ҍz쳠M�� w;"�K�[�0�X�<a߽`�!ſ��nf���;�u��=�Ej���&Q#.�+��ݛhM�s���&ۻg�ck�Go4��>��@�s�z1[��n:�T��&³�yw,[����	���}mj�Q_��ȍTB�ܬ�Y��.����*�D�jf-[���u�훟���eh{+kV��kg�Z�F{����M4p0�NY֭����s�_���.'M�퐄Y�uf@ֹ���:G���oku�lm�=^���e���{��
����
���K!q6��������]a�㋘��>|�����rs%8_L�T��]��?"H?V�+r��0�ۚ8�7�yU�L����<��0���-Ǽ�s:4���p��M��J��L+�uJ����!*�2���Y!9ڙۅ��	�V\�c����w"E�W;p$��$R����f:���AXp�ԑ엄l���v��`�������hnOD�Uq�Zq�QM��"�N1]�6�g����@���k�U|�2�;��@dZT�����8���"�1A�'��+�b���p�#u��tp��V�9�ZGdD��d&��6$w��ߨ��a�m
�>�gk-�٨ԝ����R͏j���HMe)�P`1��*&fF����i��-f0�%>�u&T���g|��(?y`N!.��D�q��F�t�����{�g��:�+ xb�1L�C��@]�6���?=��\�"s^��R�X3���r����e�QH+���UuY���yi��T�L���<^Y�M�}�=�M,0%F \d��h2KJT=�t3��E�B�Aa�LB��a$Hƞ�m��.�T!�y1̈~���M��ԮT��8�-Ʋ*%�C��n�F���{���Z$�7Ӹ�6������-�p�h�2r<d�tb�������W�����̭�LR�lu/u4���|��Bz���T�j�ʽؠ�[&�&}�c�>v��]������]]�k�h���/�C
~���a��	o����*�6���xXO����g8D#�5S�U�p�iN�k�$>>�-���aߎctr����Y�D�@�y��π���x�X�0�pJ��<J�@��u%ddd�f�l֒u4|��J�}QI��[HAM�6j1�<f@�t����P�pk�>ƭ%rub�,D�K~^����݊34v��	�o;'jv�W�v��ͳ7曬��y�&�N�����s|�-�a��u��ˣK��NW�E=D wma�����l#��l���y���������Y ��dՌJ!��^��|��~��rOB�
֠���_g4ݖW1��Rg��*S��PF�`�N�LE�u��r�4��n������"r^J�4�U0�Kk3M��=,	�R"oby�Y�Tqnjڡ�:���C��ן����g{�=p�N���u�ѿ,V��(e��O�{���bP�G��m������L���}�Z]�e�ٴ8��Mg���L<sm�-�C�{Uf[��,�Fi	�B'�CO�|,��[&�M�ȯaqԼG[���n���O�)���� CJg: 5Û٥-�>V�筙fp�m��D�n+��)i,�����J#��%�����Ξ���Er���{��p!�[�x�D;���5�c�  <�o"��6r���˨�Z�l�(h�AG�:��&=ϗ��pPe�+G�)r����
1Pߤ��噲n�^bE"�tG���EQ쩬q�K�輯0S(��ke�P"�+�f)�c��R�%}6=k����|�,I�i��'#���䖊l�Ұp�\J�_� ���^l6�LF�{���En"�
�6���(��GO@
u᠇;ʄg�,4���A�}�;�d�6���ڙ"�@Y�Z4~��a��{�i�Bo9��Nya��2�ء��w���hf�
��޴!��8�/�P�Lr��n<�eD�\,�#�͵m�{x�3�x>p��&>��^	TCջ�مwP�sbR��>��U��?_"�N����d�v�Nf<��D�vΐ����*��K��O�XUX�4�i��V3�<��顺���Aػ?���~��}�����I��Ͽ:)͓Q��-�}ff·��Ji��XΙ�KY���a'�.A�X�V�����b�6�B�y�W����垟�'��(kd��y��db&���&X���j������p+�0��T��C��F���¢�-���Oƣ�	ʆu:'z���rC���'�mg�b�)|񧿁�
Muj�}u��h����xS9k��PfL��<�E�tsSMc;���e���a�Q�沑���E�v0a84!f��ND�0X�x�.�R.m���w�3G�:�ʃ�`� C���hvWDE(����r�0O8��f���.[��W�C��i��y���M��Cʒ�D�ô�Z[��i�p��!C���f$]�i~]�ǉm"���sc��-�
 ����}�U�\$��Ij���9c|���G�����q�;����.�lwb0�E�f�qN���� =����.�Jh>�G���*��7���)�o�Wx�j����B�:탟�麘�R�eͷB��wषFz��_-��Dt���vHB�!�� ��ՏP?�	
��R�X��ZXh���$`:Hدg	0n��q��Ji hW6�GA��B2ק\I%>��A�"��T|, �^0w<#�0��[�d��-����[%���uh�J����)4E6���X�ssMe+������t?�_��P�k?��,Rw{`I�I���ߢ����q�|��l3�]
A⦎�����'��5gҸ\�0h���
9o��9p������(=�~����7Bx�e�h��ÏS�qq��Yr�y�x͕|���c>���?#����M��ʮӸ����o=m�����dH�SބO�	q>�9-W���9?��o#�ؾ�`b"`�Y?��O�?	i��7��E1� �t�u�S�f��?Y��'�_C�+�V���&��$@�c|ju�u�����؂����V����T�E�x�p!���ol�r�������\Ge ��i���eZ��6��*w5mq�C֨�4��<�3��%�Y��~$Ԟ��}���o� ���u�&���<�-T��J���	\_�~�<<�Dx/�+�z����<��d��-BOǀ�28��Z��u���(�'�ު�����-GI�eb�j�f�R��	�N�)de��Gsg(��P��j���b��%�?�"x��0,֝_ /�	��?[����m{WQ:�:@���!Q	'��� M��BR@�#�]D	�B9��C:چ|�}V ���s�!%`E��d"8��<W!�۷$�Џ�x8ozu�RDv�2���p��\����S}��x1�8UP[��y7����)��W�p�opc�4�������Ě8���%f��D�n��2o)�C��5}��R\����s�2|�_9�f7D�\/�0��9�e�v�8�P��l��_��{"�o���������e�m�`��ߵF�D��ه�R�)|%�GJ�=���ِ���`��I?䈤�X��%o^0}��Ayby��\�j�Y������Ff�O{M�]J��{�u�Oq�mO�䕦
���*)�o�8p�����2��ަO�m���P�����'(�Y����[1-\���%��y�VnA7Cdߕ1�Q�;|���7Q��=��^x��a4���n�W�	?[��3�3�U�P� -�Vb�m�\T�LQ:i�z���+����{/O��c �s�Ѭ�&��P�ۯl�ob�����/U�ʖ
��?��O)�
2L�o'	��H�q��Ҡ�wJ;,05�{���r�
���l��W�Ax�D�w�J��&&e=_�ɓp��¡c
D�Z!�o�p�����D�"(��w� )O۲�،�F��0i����h�r� �"�ڱ���f��+sR���vS�g�B,eԮ�"|7̤1P��/U?����-z1,^�I�ߞ���$a���I4�?}���8L����W�M}ɨ�,F��
��r �%��nĔ_p����=��8��"�d/��}����C�����ǣF�|� ۏ��xv�u�S&�A�����M�	&<���*FL�@�3��!��N���͎���altψ�BO��І3N>p��q:�˃]��&V�0�Se�n�a9n=�)f�����B�^�z}�-h�1p���M��
7T�\/��N����	?W��H�UƎ>����V� �,��s�JDYl��gE�p�B7�A����uը�Z)�H���&�6�$b�`ˎ���p�YH}�-�԰�j#)�%�,m�m���ޞ�
���o,zE�<�Q��t��s'�,hR<R$�ԾԻE���g��ᔋY�TkO������j�4(\M���C�6�*i(�ʭ|ZÔwLN!1jm7Y?�)V7��Ee&��DnH���%2��n�"Nͣ��帡�|��&,t�ؔ���X���۝��+xf6G�@:����78������+
�6s0"X�5�2�*V����گ� Q�~_��f�?V�&l��\`N&���.8bt���?n���z��Z�E��qW
l�2��)ӏCO�K�:�@&�T�`{<�*9�%�,�:M~dP��-�˲cc�
����l�:�B�R���^~FSʶȊ1��Tig0ͧ��w������cY�U8���'�{�5���
�5�����T��3ޟ�_ι|���5�O4G���Oj��@�x�3�)� w$,�^d7��
��V��Ȟ�U*z5c��f�=�L:f�7p6��8H��1��կ>a�cFyϪ�N�"x�"sHq�&>�1m�i@��/���kI^��WnW1�v��s��1�v�k?(z�Y��.(<6~)J�j\�kk�ܪP� �������)�::�W�E�^����t)0��Unҫ�����ި�A��l�P�y&��	�w��g� ��^� /ہn啌P�_����P��_���9G�@�S�`�l���rk$gg;>�R��A� ��M`�Ϗ����:�X�`�!��+{����EP ]S59蟾E$�!& ���M)��N��#Ws�d�o�#�=�A�z��i\�Q@IZ�q����[lBx��c�e� X�ǉ����S~��"!��iL�����ױ�U:ZJh�]��7]	����M��+��EX��l�?���n�k�:����'���A#���q��m��Z��H�q(K1܊Jb��#�p
�vb!U%A�m��n��l�֭��	be���E����m�q��˿E� ���5�&�,8�M.�3U����E��E����^\�D���I�oɷG�5�=,6м��v�w��y��-����y#�˲%f=K+�4�"�>?�ؚU!��N�ͮ�	�,��{8S�~{,}��iH!���3k ����!��)���59������F��\���h� �Dm���nl(h�"�������xr��hPBC���~f��8��/�e�f�͵�X��[촭�JU��)�a���Ʉv�3���(>>����ƒ�H؆�2�")P���Sm9� $���ř�ƴ��q[w?5�Qϕ���E̸�	���;�@�{̰��w\�	�?�������Sow�2��T�,)����k����C��������Nu!X[ȕ����g*构�0H���c�)pNqA*�sCO�K8�k���]��hk��?w��C���t�f��L��'��Y���cw������~'�q&yd:P����m�Z�����7�`c�<63�m���9A�Eè� [c�l4����	��8G=�|�X�p�E��͇��Q-)|X)I���V�$i��D�ج]���ۊ_۬�C_�풯q�~�[�0
�
���L Y�R�.�Q�uCoj�'l�cl<mn!�(�'�:�y����/E�d�=;������΃�
�(*m�sR������O��U���'�wd��	���d&�EU��<C��*�V�5�u��h��o�Q�^�х~�B�gh����:P�x`�(�D�d�W4�r�GN�����t�d{�#6�j����j�i�)����!�����hh'k�'�N���i�[��������O��N3�*e2�Us���o`AVl�GV2�Z���{-�Q�T|m9��B����T�89��O!E��;h�������D�6�9�9���	/�6����7�'��4�R2'я9�}4���5/�&'�8 �/���8W;���i�_NM+k���Q��!�[��A�ٙO?��F9��Mm��	;��"���my�anB��H�٫���eڛ��m��B(�RY����<Č�o4�oBwKgU��j��"_eFg��"'�6�t�D���X�QhU������k�#�~��u$��W���j`�/���� ���v� }a���1�����$E
���񇮯9����V�]fGI+��C�{���9���|�B���l�垣K�T���k����ϷtT�d2��s=v��a�c%M+P6|�i�-p�v5��>lzi�K!�*��坪'Nv�� �m���g�L��0��p�>z�@n+9�j����u�Bb���X�EG=�Bj����䊁ޑ��]&�e"���ca8�:��#��P�Py�dq�۹�j��h':	�Hŋ���	&*�d$�\�
��75#%&��Gp+6�0�U�aW�g�	,	�c$�� P��TK�=e�q� �B8{u����?8�r<V�~@�����>�1�aH;c���E�kш�Z,|;����6U�^�6ZA~r[gKst�oMڦ�k��u���ЩNk��5��e�`��zv}'��-�ě��e�ܸ%o�v���*�o*���Ď��E7v��%��)��9�v�ߦ����˂�V�_���7d'3�F��[:��3O��|�)���-OͰ�j�u�V�k�?	��*�I<��_9�ٗ�4��e׎�.ٛ>���HԲPβ������g�I� h�>�x�HF�B�T=_�|�G�g�m��5�əj�y��_�+A�I�f�j�Adh9K��{���M"?��ctT�����yV�e>\2�y�QMˠ��4���b5c��US`	!�٠�a!��#��CS}`�C���|�|�� ��?x/Kc�r#(�&���;N�GU�:UwO�=��*d+�a��
��\�ɳ�GQ���'�W�D�� �Ȕ�9P�h�]�s����pW��a�qI5(���fiZB���Ў�s��~5'T�s��:o[H� %�uw�{s��BU%L����Q���lcS���3U���-3�^���c��&L���k�ɷk�P���W�[��s�}�7�˭���m�tH�5�;��8{��ɋe~�+d^�Ɇsg�">�zu����l��M��֦gֱ`�ב���Yfީ�iЪ�p0�Dew<���:L'����1|Ł�F-ژ}ܯ���'�E�W�r�Z�zn����,�	j���,�1��]G�����Г'�1>�5�9�BU4�����7;8	���]X�!����I�V��o����~��ЈM��Q�O�;�`oGI}�	+�N�!�h���A��c����,thi���&r��'2o�=H�yH/���}���8�=�X��Ƿ@��n����M�`T���ٹs��ռa��^�����#sS	���MX�MS��Se��Z��>���}D��#LNOupuq;�#�y�����A��Gs�-M֛����͢6�w"��Ip&�UªłU/9�O�JZM'Dy�dL��g;�C"���@��>G��ҩ��!��
���R��S<�7�2���]�.�o�o�R]R�M�Qr��u���r�ЧN��!�ݹ������T��deu�$�$�5�z�
i��{}}Ӵ�{DG��rmQ>���-͑�߁����l�4�O<oJ��t��a9�֔{�K��z�H:�vֲI�����l&ztX����۷%θ���V�����G�!��R�1������݄����W�6��|�1�%ٲޕ+�*��6Bm��`)�o�y��?��
_�:=lf|Q�~|�����E�ߜ��Ƅ����S�Ь3g_�_z	����9&� Aoj�]��R%djU͌��EA��9E^��i5���%))�DA���'�(������Js���_�8�ST�/S��t|�]���h�lg��lٝ�1L�Wu#��'p�I�Ԭe������g����Z�qr������|����>@����ѩ���n
#q	"�[$2& ��m��)QV_;v�븏�G� ��\���'yp=���C�/�Y�e�
5��C'�zq��X�֪zn+�1+E�|}�7�U{$r���K�46<��'�|�y;���v��e��~��Hݒ�K�p�" `�>��x��yт���9�]��vyR�����˞c�m,P Ӫs�-)��N�#���+�+�u��sށM!��R��-j�����޼kB�ݐ?�i��|e�'��Cm_3���U�(m��&lEI
�I�b��<ƲB$9%1�|�k�U�QfF��x PX�q��X�޺ǵS�����ԧ�����em�+�i��+�9��F������&Fޔ���ײ&��Cn0������:�)�/��{�B̥4v�����NI��U�cG��L������-�T�ݿ��|ބ�l���@%�ź�/��︺Q��L|򡄹Ε�H�[�R��\�c��1��}Z��_}fQe�k7�� ,J�Q+!�ٸ>O�,����>�Վ�o�8"���hwۄ�>鏳��7�Ӂ԰��p]7r�� ���&f�ʥe���;���6�ۚy�O<R�'�-w �~�����A�G�-�3�$ln���.����NT�&ZIg~�����r��EI>�P�jWQؠ�ɟ�?��L�~����\ad)H�|{��9�-E�s�� MŴY���_^�,�ʴ��AP�'�� ���8�{<��O�R�e���#>:��2���*���!)v�&�Ll� ,\�Lw
�w�?����S��X]C�XV��}���k�sG8�rb�\�nq��m1�� ����®X>�k�Z�l}�`
�'�S|9�����j��Z��I��l�����҄�}�ggdE<�{���y ���|Z�L��O;X�������Ks���@{���:�E�:N� ��=�6�ȟ��0ɬ�����AXg�֩��"=d��� ����szP9�-���\�:�DWPĴ���ף3���ʭ�1�k�+��h5�k�/��³��̵)�:�XPd�U8�۬�� ��5.��)|���}�m�E�1��O�"��>��d�ȣa?OKĜ�7v���eA7�y�3Ȱ_ؐ����gUҢ8&Y�{d��.��m�lΤPG0�Gl�|d�����*��cUZ{����A|
��f/K����G
<����a���޻�)�?�9��4�3wa �Qb�N0v}�����}0E0B�EQԔ�QCt���E�ir��K�טD��$�QG�\��
f3i��tD�k���7�I��eE6�F$2٪ �� }������ӌZj�p(H�E8�����fh �W��Ȱ�r������a�#1�����4M�r-&J��h;�̘�W���VΨ�������������&���A�X�A>���j[[j��_|c� %�͜��X��j8���1>�n�]n�:�MK�z$X�*�2r�3#�� ���68�z������Q�](r-�C9�����̽=
t�-��T�f��A�����>�[��|�$IZ[����b�v�p~��RK�f6(�0xɏy����Ǹ*[�����3;�|{�_��d$����}�p0�	SLP\�,�Ƒs��YA�vU��Y/�t;���ܰ�M�V���i��ԏz+���K�{��|%k�d%��x]��}p���R�ْ�[ne1��1�F��
(�_A!p���F2i�xެQ����'c�Sb[�gP=DӉ���1�/�| QqF��W[�y;� 3-8ѷq��ö��NCt[�QM����̌&8��-S��h������O�Ф(�358!��J�BF�kA���=��{癀U�[`j��](�F3t{�TYK",�!I���O�|�Ơ+F�u`0���SA���B�Tv���|�(��(�M�?����dn��&w��L���nхl�"m2��hɥ�I���pdT8���nӶH�Cr)�X��w|�#7�Rt�vA�(��L�4
;��;X"b�PRyT'�^Ϝ���S�����zҕ�@���#�U�,�&������m_�����
l��Ò��{���c��y���H���`rr.�x'�+U[�t|�[g��U�F��;r%��'��� E�SLd|�V[i�#�/��W	1}.&DT:����M�&���!(I<�z���d��.j^N6ݞT�����w�^��Mmg�����w�Pۃ���#�#�b�s߶�l����p��/8 htz�Нor:'_�w[EpAљ3��h5�
:�
�z�ϫ}�F�9Ӹݬ�O�-f�}����d��nS���bW����:Pl�`+C�i�Pz6"��\c����}Ak+eM����h'�#o������E��~�a:kpc_M�]A:�)�$������o�ʅ>BRL�0�Ɩ�!�7�J��}�BdK{SX5�����vt�FV��}H��=�-(&�:���F���b��|�1����v�A�$�X�����_h��;�s/�	���}�*��_�K�[fa ��M8%5�̏J�����R�ׅ%�X$Lw�I:P�xn�<��WU��Z?�Q ���3�PiH�;��X��P�r�ɥ�k������LũY̻uK��>�k�\��毢1s�0I���Џ��w.5�n��`w�
	#�֨�@P>xNk��*�L�h �:k����k"#S�.�;�W�.�雐�wL���u���R*&k��� }V��p�_(l:�����؂�I��#=�;��RX�b�~k���0��5��I|ʖQ�θ�u��6@�a3X�@�4�A����'�֬��:��M�j���>�''�����c�YTzܠwf�jݱ_p�N��4H�whf��o)S�Oþ�p�x�=���S��Q��e$��S���+�3ٖ3h�h�\�Ͷ��݌:�`��5h�Bk�x-ף��L�f�"8ݝ�	�5p��������
��J�&��}g���Jm�����3D�1l]�O�����~M��\\�����6 _�n��tHc���܄�����

8��\ � Ž�v�v �PG*��o�[[�򟗌�V�����k��n�
a�T��ɰ�=g@n [6�YP1o�ũ7����f�k�cġ����?Ѻ�M���X+ԯ����e�(xDJ�cz�[ctK�u������X9v�ցsq��^��[d�����N�U��#��ѥ$VKP5�"'ז�\���	Ϭe��̛��k_��¿}� 7vF$�g�?x%�M���$��H�c�[ՙ���*Vh��,�Ǔn�e*u;�>|��,�heG#��A!\���Ϩ��)o����5Ԏ�]�;!E�oL�FE��+bM֦h��>���i�8�N��.����&]�j�6�O������k2}J-#�w��زԿ�!˹���~ �����c�b"��]J�e�^u�����T;D�I� \Y��$��6��-N�jGmѐedFjJ�	-�*�򻣡�w�:�� ��%�HQZFQ"��<ے��͔�"j��c�#1������V��^Oo�H(��r�/viϢp�b#u�**�`��+�d2.���d֓'c*�q�/���H8�0��L|�]nCj\@�V5&����G�����e�2����%�&C����y��">^�p�r7��\�3���̛�u�W. �����=��\d3=���u$�OSV��WS�^���0���!��ƥ���rL�_xk�8�
$1e�Քr�
�e��] /Z}ܴ���
3������Ĝ�#2�ĥ����U�M��`��^����\b�n�p�4ݼ�Y�#�[�9	?���8xQ�FC��������j�V�I.����>w�n7JuNC���.���`��b������lz���۱Y��͓���3��?���,�ɜg� ����A�6���������G�'�Qa����.��$� 5�):�����FN84�%CiR6e}0��_��]�QʫYؾ}�J�7�"�9���0<���o��h\^@��HI��Űt yuߋp�����|đ���K��}#=�?��1�C
���ͪM�e걉��.����7��X%,_�"�F���>�g�B�;*Ұ@�|��
&g��\A�U�ӱ�x����'d�-B�r���G0��*���&����	����jEY�ۣچԺ���4f���`hk<�[8����L ���	��S���µh�K&3��.�I��hj|����6\m��#�;�_<�����]d��Wu��	��������^�5��2sr��L��-� �O�g��=�C{�H��
��3\C��s��0������
�.�%e�YZ|�1c#�ռaeW�T�)�:�CB��EG���_خ�	�ǁ��#�n���{*����aʵ�I"w���m��j;@����U��=�Y���&��
��Y�c��[���9��bp����PM-)�\(�\��v?MSXB�o4�Z��F���b-���lI�+�n����Q�^*��C���;Z,��B����mo�/�,K���ی~����q�
��E�ea�������&+9�yH\���X�X�Mç ��|y�z�rI�*ذ�@���zѭ���A=A�c�=�k�P���4['�R����ܸ�y7���ֽ��4UՈ=E�j���5Ag����t9,r6
7�fV��8���`岺.6��������Wک�6�� �[��#���]���v��7�����L��`���.2*m����ԨQ@�w���k��E�6�w��'S�g�c�����:{˅�-���W=���wVA�_
�8+�M]h[��.� h�[���b���ܬ�|�}���'5��}+Fk���$�9�V���i��ZV�ĶI<CSb�����R*�QU�t�RV���UZ\&����p���^^6eA��n(��^\����h2#��������O'rK^������dC������9B�6�#0Ӧ��)ޝ?��ڒ�\u��O�_��T�x��CC��
Izrx�`�_B�K��
�㭋��)+�� �`ܝQ}�[��ŝ0?������BoF/U,Ր����f'c3�����+�0�sC�X����鄕J~�B%����tv���d{Vy�����7f���E��j��O�`&�"��D._5��e�"�ޤ�����������ʠ�� Oj��VzkA�b
�'b�|� �8U��%��̣��)a�y�[R��~E
p�y����1��ɛ���M����wٜrOd=�Xk�u)ZJ���JR����b�Lx@���{�	�`�7'#��cE�
XR�Ll\c֫��m����'Ǒ��0��A���#>hF\�ĉ1�!�@>���Pylũ�K�$�{ R_�U'���	��ۺ���@D�\�0�W��bgĉ��|��Xr�!�}=��.��� �H1�Y20V<�0���lPmy@����P��{��DܺW�d��L�[���������+�I(��捬V:$��q��Q�A����q��߁�d���m��v�qT�sD�Q������h	a�DG��C�Z$RK�`�Me�V���<���p�ym
�o��a{�绌�\h+[p�"$��0��kYq��e)�v�%"�7���sDn��)FD��Px ��8nK#ѯ����g�ǀ���>�$�]�JXN?��2���F?��4�_BX��o�ܴ��K�b:�u��BVb}�\�g��)�e���C�:�{m����'��䰘=;����ƩMQ��%�[�n���\F��%��>z��vuc���?�����`cm�4a<:'��������9��ҏ�~+|�����c��.�=�v�d����Ѓ.�,�Z~(	�s��q]�np����K"�hƽE%��7OӬ��晳��ߣ�`�����%�uD�"Mw��p6�8�����O�d	)u�-*��H�4�s���c�t��~�cuP�(��9z�L�{�#�-�6P�a��ª<�q��6��k��ɐ�����:�d�lR;��\7�
ס��&���T7hUgm��00+��v�m:�P�/��҃V�9����/������"q�}�rW2�W�B �AB��m�J0\�(vj.���Y	�F���C�J!�Z�M�d,G�c^S�F%ؕ����`�u�}2Bx�tp�'䬋PQn��"?�>���&�$�ߜ�V4oI����{�+^����ti�.N]�?M�i�c����i��мHe��B�5�If���|��d/ȽRܯd�0�b�(n�lwkx�8�����+^-����"�w߽� {���>�2
<�Έ4_?f矩&M����8j�g��w2�c z#�='�d� ��X��ε)��q%�Y>.��(���w�m*��r$*�Z�j4pDuNk�L��\����/�IjxTe��x�� &��R�x�0��RتY�Z'������  x���ұu)�PQ���_��t,Й\�W��9%��jߒ��BbX�Ϣw���`�͉3u�(C�������֒K[�p7��*h�k�S��x#<Ppf���	�jR'��@&n��z��>�o�s'&�N�4\�"��r-�7W'[b��}�*�axh̆ty�L��Q��>���&�n���"�/��jOIsէ�q��ֈ�⟴��/@V�h����/�J�}�в�x��m��Et�{9�`zM�`hy�F=��Ҋ^�-�}e/�[��7�659�6��{�aK�Z�z���Օx�;�TBd�S�`�70��}p����yO�T����ʌn�03��:���13K}W�W�u9mQ�	���qu͑Wr�x����
3�f�hw�GmM�J����ߔ`�Š�$w��K'��nc_��%�!�a�^;�t(�Tb+�֟WW洅��I�)��V{��,�L~vA�G�����7�����Q���p��:���z���[-6�g}L��ō��Х!-�VT$6c|A���#��D�1$4'_��	i6{QZ��-�V���7�s)K�N�"�EouGs	���?�d�2-��H����T��<bЬ�s�:��7�8��!��u� ���k>�B_��=ʼ�����Z�����01 �LVIO�|N3���w2�8#�!�6 +��&�;���Т@3F�χEx���|��,��B�I�t-����?iۀ�m�,?���$%�:a����L�EY{lc�)�W���d~��bߌ
&�ۮZhS�/	Sì!~���^�z��#�Hd[y{ҳ������.)w�O����l̃�nM2�t��]�����Cܦ0g�����o%gS�mB3�ڄ*#2f	!�+u�|���K9�h�iI�c�V�6�N���=`,�h�G�f5c���]��ڣ�4#��$9��˶!��0�by��Qr8%X��S�2�����ݞ5>��ʚq�n�~B�ہ<�,�D̕���W q<XF���9N/�ˎ�">%<��,5�Q
4~�sz�塮o�5Ə�8��9~�h}[��JO����r߀�pQ9��!�Ͼ_}����/�K2�]dhs-�%I������6��07��(Ъ�!<�����*�ʼ��Y�u�
5 �Ah_R~���BL	�Q�Ƣ��W;���� 3\V>��=�_L�JϬ�d!���}0f���P/W'jz�5��#�5����` 4,ď�P��nN���%��L�t�3��A6�7�x��`2���.�>T]�Os�<��Y'qg����@��1�9�9�r�)����A�z����t^�4�d�G.��_�ùb3)��Ceݏ�Y���c���c>d��'��>���צ�&�˧��W��.����ӧ\���*�)�~yt��
�� j�������fO�⧹2�z�9�I�4F]�b9(�m^����^	�nw�Ǹ.�{�PhLn�w����>�il�g槠��Z��΀�"�g��(іk�9��n�tM�'�Ƕ����
�w?��[`����3�l��𣛚^#���x��$d�.@WU	Ն�E��<��ɻ�R)�H�[�o��-z s���*$��jvk.�6�l�6���o������!��7���w���n��A�U��P�=�y�!�&`�X����Ya�����V Xeb�;�3�}��)ۤ+Bج�^%�"0)��8*�*Ϟ���a�������AU��߸f�e��ZhW���ܖ�IB�:�Tߨ�(-�I�=p@��7��h\�'�Y�E!�t��¿�K��i���Ea�P.��0ֱ��m����-����=Z`A����vǺ�\f��l�zv��t1Ӿp���n8�ٰ�\j|BL4Eں{�>< ^���<�Jp�E��:�?�d#�t��JLgw�7�J@Q��v%�{Vf�(���<���a;pK���7Tψ+&��F�@���(���dTv��c}	A]w�Fp�9��dMp��k��`Tw�V��&���|u<X�3�֨1�� �_�����$�����$�P�;V��+N�bRz��4��̖q�>|�A�������=|�NZ����犚�6���&̀$a��a�~�y�����IZ�@�qb#!I������J�d�} λ�/�,���Y�i^�Z�<��A6*�=�2Q�7�䡂s��x��P3E��� ������>g�hp��)[)�9�C�^ ,'d3��e��Cj9�ᙯ⾚�Q���{l�h�]��\��Iى$�۸OwX��
d���x�B���w��a!��Q� �E���m�J4��	ΆHbd���:F�E����VV)!Y$/Aw���`v�M�7wH}��gN�4aT0Jq�X{��9e&�+95�XY竳�"��c$�nm�?���������󿪆�eW��G�@,�ߦ墁�8�Xr�Ix��}CJdt'��F%Ba������;�޶�~�r��J[b 96�LPW� �m;�}�
� �Ҽ���F	8���@y�g�ވԳ{x/��2��R;�T��lTf����p�:���^�0���Q��v�9��%]0�HՇq@_9t��h_Y�I�{�Z+��Ǳ�dXt�E��"��0��j��<���X��Q���G���PS�Z�f.T}��4HV�5��4�zQ`(����z5g�7=���,��q2��8�3��ctg�Pa2>�_�g��R��l��
�0*��Y�&���u��&��o9��V��K�������`V	ܕ��}V����v,/ά����u�� ���I
o�e\Z�+)���a�R��M'�{��<u)[�R��\��B*(��X���Dϓ+r|�*�=�Y�;��z"���C��4/�FDс4�W�S�����;�& �O��c��u�Q��H��e�%�Yh\�Dpx�K	 V|ƴK��M���8\ �������؄r*ەǡ�-g~�ꔎ��x$�5�Ԏa�^h9�pP�������$�SC�8��:sr��g���s� ɑP��Z�d3aUs�[l�M��1�"ċ9�7��o���r��!Az����������'�����bZ��U��P����nN��|O����O�C�Fo�p�CcԨ���^�4=�J��|Jvf��O������gy]P�#y�i�\�t���s�oar�*�i!��!���1 �(O] i���f��@c��Q�M�_��Wh��LZ��?UJ�O4��LoyQ�c�����I�8h��"�Z�������6�i��&�07�D��=�lB?�Л�-6|M<�/�Wᶡ2�z�q�mg 68��	�F�����'ّB�g���r+�{���2�°4��Q	����nB�c6+=�0�"�VmYM�ڤ�6��J�7�b�wd���o�i�0�����j�V�4�]ْ�e�]��I�էP�|}���s�leddO�������
�*7�.�6F�8��j�+)4���C	�#Y���M�.D������p��<�:�ʷ*�t�|����NDL4V�Mz��R�y��O$���<�O���)M�xӃ��rȻ\�,p���c��eLV�7�Ңj�Zԃ˷���·K�.�4e�V��;P)�P��|S� ��F�^��K�͑���x��s�(R�a�x��h�t�����*���8�!���l�rH�����X�G��p��1Sq�	��.�~�i��}9 ,j����Eo�����Md�C�ɬ�~�%Sb`F�Fm���tc�F�a_M6�,᥅� ��Q��[��˿/�qn��>w��ª���`@
3"LK٧�$��<o�cs�T�+Ʋ���s�Qx�}'��µ�}��FU�<9���|0�g\ݽL�s�����e�����"�Gw��|����n�V�Īh�e���y�O�h�ŋN�;U:+˫ ��D
]�e=Y��G���w�8���������r����&Q'�ݝf@�Ƚ���>E�� Hy�Y�r�"6qJ��άYE�}�Y���&��js�:�%���ig	/�H���s�9ř�}FL�ʼFKmR����H��ߩ����T�v���N5;�4���X%2�F��<ҵ�}2��cCa������KAEH@�*jT��> ���}�TTacޕ9���_����>�����e�yk�,n���ݲwfh
���_��?Ui��~��)��N~ P�/A���~&��d
,��BF%k_�����S�TH���'A8���_(�i�c��Ė"2��˘N��u�\�M���0~^�"�/P�/�@[�O ! �2�%��J��PB��H[�h�Ml����9k!x@�y�b�IDU����˄�'R��;��� ��D���t��cjV��7���[J��b=�~$n+-M��ojZ�v��w�6{v�!�V���e����M� .�h�|j��	�*���m��7ч(�3Q����r��LB�%#�Lbt�L2�2�W^3z�^\Vȷ#M�����H�X��������p�:˾�|��:�������B��?O�.+!��V��a��O	u}{?�P�z�+��.��8��^Mu����� `����V-H/5[�@�g�����ag��5<�SS��}������Y	�s��Q����{P�1������&+�c�֕�~KR*UQ�yi��dױCq]����h�����kU�m�#D�^�*��=}�r�
E��F�&��m)�q����Z���o��\SZ� L���A�@'{�?�9㡑|�f3�os�VF[���,өſ���_S.z�%EA��au��B�k���\əf�N���?�Į�݋W�ߚaM��8���{��ߢ��ŰVa���[`w�d/]������~� ��O�f���k��|j�?d[M��l-HU?�{��p:ǌc���,1���D�V(Ps��ך�1��Ua���� 8xV��!5s��ڴWN��|vV���~0X�<���)�֠a�\�K�o�cz�����X�#_f�`Jc���h1cH(gį��fl�'�i���Q1�����C�?���q��e�Д蝪=�hhp$ad(o�;v&Wv2�V9aqF |�Q������綮Z�������7�;��y��j���0�2B��5����_�ds���?���/6C}]	�?I�d�s]���X�#ᜥG�e�7 �SU�<�����*�j�3S�3k�`��@wK�Ymj6CJ��2��-�[����w�'	�Y~�a騷<��̚#��$tS�������9�jl3�	�ZӻQ�#?�/'��TR��x��LW��V3�;��g�hs��7⏌�#���	bko��/�eA
��n�	���J~�|n�aă�{�Pג�GɄȾ�n��x�#?^_v�a"��]9���UQ�HEGff��c"�k����)t`,���g�07�7�?tֺ�e�$˅Q�l�5mEV��00f�K�RoB �)?��Lm��7����D刻�Þ��5�R���p����5�������$�F���۰���E8I�먻a:��f�+��W�5pG)
2��T�v>���9^���A�vľ�q��!�3c�>l��=`iF���=��Is�Tj�`���i ��/���R5��.��=�;��ݺ#�#Rm�?Y�ч;r��{��54!� v�; ,=`�$}�Kz���3�Y٦��q��0,�'��s��,��#2��i���Z�D��J�؃�{!�����]����@��	1}�'�>Hgg4�ҽl��#��{���KeGOLbw+G��PR����0�O�
�f?�ٱ�x�F�M!Z�I�1,��0ě�*���*���Gl2E�h�8C-�B5���4<@F�H�X�cf�-[��!�����Ǜg�*NO�{kW�o2Գb[�!�v��2n�MO��G��a9~B�85ۨ���9�����N���k���NB�t�M�����Ų������+�fLwo��\�/�v�u	�Q�i���Շ?(�%�R�[#t�T��n�'��5��.��M�:�ˋ��+
h2��Ɠv�N3��	ĭ�I�����/�W��
G��/���E��P'��X�+�r�/�nZ���p�/6wY�V'˨qʎr������ȥ���}�������2V^v���-ą;�n�z����CՍ�x��b��={�A(q�*} o+_q� B�{�� (��f�c!��tB�SL����@J�GxꉕfM��?Ƙz�:>��!y�%�}M�{�Zh�n��F����d���s�z4
�3J��|��
/���|�o[�F;�n���_СyP<\i�ah$�ާ��L��֍* d�]�Nk(�}�Yx��%��D�M뵿���]�w�*��Mr�����D2ɃIWv�j^j�^�	킒�-��5u�<�e"�~���e�a0%"��KK!v�MM.���l��%N����>=N���?����7?�H��'��zR���\�:�nPY0Q�p��Y�N��bD&��5��*�8�4��W͆��%RW#�ޟ�>:���8�}�C_�=� �l�)O"j^�ʤ�@�E�aG4��IY�U��ޞ�cF��s��U�^:���J�A�����F!����̛l"��̿6�q2���d�/�)��^Z÷�^y+Z��3��RQ+��eDx�{'=8Dա"�k{:�vM���S1�u�K+��'vd��>,˔6!��1�-�r�qvz�h'�mk���9��^BW����zx���G�O�۳Nj�%�Y��t�q���
��Q�Lޣ�Ҹ�I�.пR�����e�e�h%��� ���5uЪ#`��V��L۠�X�O��A��Soy�������肋�n�0��+0���+@j�š�l��' 
��6Ԥj�;Г~�ϴ��b��dcX�ǽ�����5*�v�pŖK�M�����׼�z����*�d|�O�En��)'��_�nFJ ʺ�}��PZQ�Y�F)V~����Kͻ�4����ѱYX|��2���b\�<z�-L�3F.f������?ϟ�n<�5�����kT�b���m�_���0Ͽ�s���I8��E�4#y���c}w��vȗ�3r�z�������BN��Mj��x����-�Һg����qb��uv~l�a)ێ�H�\"2��E��s6�Г��'x�����n�CPң��<��M�"gA�g6->�>?,�[���I����x/����1	���@w'f�}EM�k��od�]�Xc�.�
�jţ���U�Ƃ�:I/d��!Q�*�ã��tRe�$~�-��0�4�8�V�/vt~��00ew)G`_��CU�����a���h\�
��u���)�g�g�NV͟���s)j�"��)Wi������iP[��ɋ{L��Q�lsW��* ��,c
�m���Wk���L7�~�l�=]�f�~�[���#�5�T]`:��}2�d&�B�"{]��"���Q�*������o}��уw���kn�<���;O)`,+xx��l��W ��6AsgAL �!s䚲���nzKw1�F$�}���X��r���r0;j�>y�F=FZ�O�ėE��8�Ҝk.Ɏ�+�p����G.�޷��O�mw���7I焆v�͏
'�AkPBn�I{�@��j3�(MA�R���7��>�$%�OM'<yS�*�}ޒlx8��z�� �w���g��rE�?k6ҟ����&���q��
m��������X�AS/%���F_i����n��<7�4��w.�lP�Ӣ�H���~�R��aq4�˪S��3��s�<� 
�lXg��b�E�+͸p�F�&r��n�'}��X�,�Q)m@qJhA�ous�Xw�=m�4������U���[���F�B.�O��%�	�EޯoH���*�"�d؛�&>���Q/���m����Q<�Q�Ӝ�\r���3Z�l�O�V�����FEE�{�Һ
]Y���۸���Dؑ�K`��Ϣ��$"7����t�&���5�A�U/%��NO��[�q9]�kWR�ݩ��\S�u��)W�C�����ɾ�c2F���ei¨�QT#�Ә�����t»�¿.j��qw̨0��"x^�*e�My/u����x�艍w�4pU���t�ݏ�mu���~@F�M���W�q�_W�lj�E�}�f#�R����=Ά5����O0��#FF��e�#1��{k,�G T����-G<�S�����~����Z(�2Vc�"9H=��S}VS0��Jlm[hb8��隗2��τ���1�#	QŢ*�#js�����x<�̆o'��^!�Y!����z}iٰ�'cƮd��~�{5�к���I%�;ĳ?�Y"������d�maBg?41D�)*y5AhЉ���?�`�#��Y�+�j��b���a�+Yq�.�{C0.#�ՎNb��S�L���
h�De��f	�+ *}����G��-��f�gDU4��<-l�X4y��3�q�4r�(����*�oL�j�Gq|����w8�4�{qYz���Ͼ(@d8��R��ZQ���r��]h��X��p�Z���5��Eb���\�/�jc�x��<xj��BW4hU��{恃�月�,I��'LyȠ���D�Vu�#�3�~i��#�<_��_��Z;���GRhMeG���ap1ķ�I������y9����Rr\3�,��C�C�}�"��E=r�Kޕݙ�/���dq�1�3��ݡ-���h��+��b׻�7ޠ���M-�3����k]�}i�w/������Ÿc�	9T��ۍ�)��գ�Դ �����fQ7:`q��c!,�d~ �d�Y��q�>�σ�/5Fg�v��������2���#v5��VA�u_-����[h�~~�챰m�RA��h�Ca�ޤ��;���<���p����!�{Wmt�?Q���1`�4'�2�}g4sPI_��8�Κ�'��zw���H柵��Ӡ`{L£�S�����r�FX�0�]�S� x�)P�2����,�S0�����v�ئ=�K0N�QW��W'�Fe�fF�_q6�!^���^���|F� �e4e����0YN B��)�.�y�"Y^����
��|��uahI�iƪ�	tZe�,/�F��s�L�|V~N��!C$�w�T%�-�O��_;�#�ƞ�P���l�?g���Y�\S�j�����=hpT�@�N�h^��Eoؤ]�6w^(�@PDz���r^�w��\oC�J�w6p'|ɣ�%T{	f�J]<���{	����!�
���h���np+e��|��	���xt�nE����;��VE�S�5�P	ʾ� �ެ��j�g�-��z��'\'5"\f��+�f� 3��^5�B�=����P����,�.3zy����������:�̏'��N~P5�q�ɞu�y��>�C)\�������y���g������Ȏ���`�������p��V�t��!<��d��X#�5݁��z��_]�H�s����c8���N9�]�"��k��͕���Aݝ�p�$[b9n ��u�'>k��UE#�X�g��!�'=<o��ǂH�=��C�(̾1+д�	u�?��1r�[�n�V)���nگ�(~ŭj~�3C��.�%f�`��r��Y]�!�nP�oi��Vد�� 	�Nʊ9�J�_�1,�A.
�� ���#A�խxgi@���r}�h�l �K�4N6���(˱J�UJ.�;�Λ���|KX7U��$�s7�l��/'_V��f��A��p�5��T�0�\$���нԃ����IT7�y��������#=��Z{+u��`�pr����������n�)�Cઠ��k��܌�3��Y���mxkO&�ވ}�����b�/qG�i�h�G�zN7uP�L�l���7�$��W>�'� ��X�z�j�:�^߼I;��D2����2�ˉ+�R;6A������/�+� Ӯ���i$Z�8r���ՠ��"�����Vkv3�z;���-��o��t������'�Z�#�]W
$>D8�c��v�[��'#�j>Sց��5�_�d�F]���4T�#_)�͵����۲
� ���4_�d�9�x�a�}��Z�-ȑt��0����$����"�㒌^�J��r���Z	�@~�4�/�,�O���{��}U�����V�e|�A��
l�U��^}[�b�d��$�6=iIC��iu����~�X2mQ�_��TO�]��f)�TZ�Æ�	.RD|�֊Ka����XJZ�a�xd;Pv�k�)�%��4�Uw�6�nRt%�r�m4Q l�t> {-�*�o�b��KE�TmL�^)�
0�m]Ĝ0<�I���;�h�v����=�@��縳�As�Ս���M[So��Պݱ9Qg�G��W�4n��YA�G�ZC�%L�R�;�»喎�'�X5�bo��[�� ,�X8�,ˊ��������E��!dKB�a��Fpa$鴿��qo��.���	�g;��ه�.A��kI<ޟvx���' ~�Lh Wy�R��=뗪��i*OMi�,�X��{�ou�i�����>��|Ӳ�t'9�������_dEl-�ٍb�朏�HȀ���WO�K��$�m�S��]�008`
6I�_��ܶ ���%i�s��&ᰘ�Kp밞�J����(C�QGD<4� B�b��Bp�<�n祵z���"��)��0����d��U�vJ��plCQq/��Ē	����% M��J�A���I�t�8E��ІdЪ�Q���0�H(��?��H�Yo���W��lq�����]�4��߆�]Pq-��7X��s�SR�~ޖ�(�Y�X���l^^����� E���,������+���9@��~��=��WZ��o�^b�J����د���l4���0��d_���� 7	��LW���4,�~��'�V�!���
/������&��7p ZЅQ4��b�]���X<�A���������q�Gm)����	E��y����+T�E���r��5mZ��牁M�!�E���0�)X�����ԃ��\<�XI��a��������k�It��/�X�A#Ո��h��/��ԅ<X��΢ٜ�l�#��h�	��@J^�d�S��:����>�\_*�C� &����i&V��Ŝ��t��$<I缅~�/��%��۴@+U7��ǥ2�4�4-ֱи{rg	T,�U\`�66��3c�LK��4����,�@a�l���\C:�m�	>A��
�H���5���{Y���}�(n�U��tRz"�[L������2�t���xE�j��6�d����/�$�"2\���$�X->�?k�⺙v����I�����<�iªӽM�}_:t������z��+-BBY��M8� ��`P�e���3|��_*0�^9|R/8ݡD�2��u�V.�0'�1��ɷV���'ySm{��VC��|	��qQ[��e����I�<3�圉Cy{�� -�\Y��E�\��<=,���AC�b�s*���M�Q��z Ti����2h@!������41x.z���	�W��e���U���U8@��>�(pk��3v�núsp�}�0ZA[Wo�y��y�7
��1P�<]��O������6&zp�^T ��)~ׯ�V�����uE㴴|�_�U��.�C���ٕ0� ��h��k��������I-�G~�Y�_7?�f��n�i�An�ueS�?L�����A��%(�@Y�I�Ot����F"$Hg���)��*i�����%��(�tT"��\��<es{�'�����&�P#0t�<����n�������U�"��
�2����t��uu�-����zB�0lƒ@�3��ϓ�7��מ���+�$��h�� ����.+Kl�x�xV��v���	�ؤ��1<b��Da!�3[�J�{�_��Bv�F�o����`����|�q*bڇv�/��&
��X��eŒ:��x㧶�K������m-	�߫Ƅp�dGIR%�Ҿrٙţ�Ǭ��+N��ڱ�(�?���=�!���1�Y�,�e[��-��Ro�'�o�D��F��/�8�F�:@��h�c�Ke@T]�r�����Q:z��8�#��#	tT��8�,�<�Ì6f4�LMr�yPK.r�0&�Nj��t���v��~��֬�-�:��R3K']��v�a���$��ZS�K�jBY��}��N���E]|`��F&R+�K�ҮB�h��5ݷAJJ[��-YQ|y��cW�$&�te<�2*꫓����>�X��p�B-��M�~@p�Pm7������ō���Ё&`OR�<�A'@Ì��ӹAee4%��P��ڋy9����^�Bs����Gԗ4�\2| �$��V �q�N|)�\��z[����#��Y옋j&��*$�'^u9K=:qayN�T;0Y'�$3��"�M�X�I@�s��X�����噶]�L6h6}�p���Z	V<=���� �
�P�^���x.b�E�l��y� �/m���-�2�� WKu4�q��I��PΩ�Ϛ�	���V�Օ�P'	1�sn�{)�E��hK�	ҳ����H���L��S�LHh�}� �o�W�XM���j���2;��r�l�m}�::�V�LņS��zĴ�r�]V[��e��={($����%�D!ϓD��(��2�������e��E�L�1q�4�g�-��(v���"3V��V�@>n��[I�H�В���BI+\.٧�qA�M� 3�n��k��X_xef�#��׽׀� R���y���<P#_����FO�z�Qg�֋��̻��@
�SP���*����LOel���u��AB�vD#��ړ�Z�DO�DA��q:+Q�br��m�P�ѿķ����q�ӌ�M\0?Q����� �� �*7^6���fb'��N	8I��'t�t��,sѾ���F��Zo,��X�!�!�|�(�m
�	��V5���v�!4�$�N�<�d9l��%9R�b::�ܛE��<	N��#�;A~�c(p{a��~=��p�P%�y�p�U�Y�.j���P�IX0�O��j��`��y�lJ�(�nM8p.;��؟�©�}q�~�P)���xeHR�j\МT�9g+`�DƮ�%t-����:��xv.	讼R�1�,uy�90�S8�f�;�o+��N�hYq��Zk�UXU֤����p\A��Q�K�ߥ���>`�A�P��҆5��Fq4��I����5vf��� ��k���~�>rqɍ��mx���_��g!4�B�2�Z)�>�}�\�.���ۛ���ܽ�Ԧ�:�&�K��nRC�]���e%��o`>���?\�_�6�^w�E�z�0F�u���S�b%�W9~��5�t�ٙ�Q��A�Qa1����
������Ռ0A�����B���v\�.��u*@��%7��]=t:��_d^�u����O�`�M�jٙЕ�B��EH�c�Fȩg�T��:"`#EW0Q�vm���o�M0O���Z����Zr�f�Zp���򮲾E ��MbYk:����y�����x�ի-ѿ���_�m�	K`�TI��-b���,��%8���P��� '@A���罤�{��Ȅ�4h�1��xN��Ș�w6xx�������џ|���n�����d�(L`j�Z�&�HA��w@Ͽ�^��}��
�����̽�����G�V���.zv6$?��ݣ �3��f%1�Yy��O�V�\���)���+K�`/�2�B2NW�O(�E3�'r��z�������QRז5�VF���5苪�<�����o�C�~��F�T�>v���F����"k:m��
i���vɅ�_oݖ[ ��BM	4\$$1���M@<� �i��${D�Ȧ9!�M�*5��jڵNj�4#��-�e�)�퉙#�%��u{5\��Ԗ�z^z%� Fv�F�+j��9�$
����q���j#n@�x�XF٧�	H9���U.Q������M����@�ۊ�] Oۢ������;.ߢ=� 3�@��G��h�lm��]q��C��=���<���b	#���\M�[ں�`�\���t��;��ӋJ�՝����o�#�
$o�vk�g�*4�x7[0�;��i�Za7#/e!�~/�a�
�~Mt��.p3MyI���Eц�:O�~����cfT��Oa�Q�4�����r��!�@pb�^Go��$w��1L��F@ӌb~��Ef1�4?&ntl����@�5��%�a�,�	�=�*	<�֨U�1f3����Yk2��x�q����\C؜��Д�F�5c�
�ts�J=C�!a��
�k(u%w	N���ϝξe�q�VB`������ஊ8V���lxʱ�4qʢ`������Q�H�q��ݱ�e�!�>�d*�>�9����T����`�+ֵ{(���S���̗�/�Ռ{\�f�D;ɛ�#k���(�(c�TͳɎeI����� ��h�-5a�1�9�6;z�����`�*�=~���d�n�Ɩ��L�yz��?7Փu����IY[�I��vX�p:6��j)^		$[+���{�qm'�գ>3���"e(z��N0+��A@V��6#
�?=)�����;t�k8u�wB1;��I�;!,v�+�%Ν�(����7ᥜ`��"�l�+��LYn�e@{R�����>D�R���z�)(��	3���kto�u�c:�o���m"�R�Eq��z��E�.]����'��OѶBSsl�����`l��ߌ9/�}ž���������&VǛgC8�`���Mc��e��,t�f�yLc���/V^��D���>=߾
<5!�/q&�)wH�D�r6�6Q؉Mb�э4y)ŉ0"����#��
&Q�ȥ�1k^�u��Q8b�R�
P1�
j7N`�,�DE-z���Hy�ڿm��nHi?*�T	_����%��0���]Hc��`�\i�嶆�[���'�X�E�;�ٞ*"À:�&��4.
|m����/�ԏ��ey�O9���Ӏ�M��2�7�&�пI�܍���!6�֪T�[�/o��Ԓ=_j�<����T�����taG�?���A(��^����z��C��~[/�����u�w�W����S/���������q��u8�a|g��p���^�d�o~
AȦ�՞��xo/m��1�!��� ��h�7Ϡ[��ʟ�B����T�W8-HtTR��т.&ϰi�ղJ�
�$�C����z'g��gC��T7���zݏ�m2�7C�!5�h7�����B�"�������`�w�h0A���U��,���a�a#�rB�Z!�Ҕ{X�M����sM?���H�G�o˦�V�O��i�S;�H)��3�f��d��A��I`Fђua���ؾ�Fܓ.�����O���~��t|��	��n�Ա��@�����&�5�����0� /�ڈ�L���`2���y��	4c#`S��j����Qtѐ�a�i@�|p��b�z%gq���0�;l���U�$�q�/&������EҠO|���ݬ�j�["�ST��(Yu����>:�YT.���}�	N(����v#-
���)��8��O���һ�v)�)�)c�t��>2�\���W���N����W˧��:D=�g����:2i�LΊ�z����?�l��#ְ��m�_�g���x�9����O7��MJ^�p�7���<��A�د'�R�{sL��?>��,I�D��oǽ|��.ֽ��I
�)*�v��BK'��sc���2�8�"3�,���;��:Ľ���AY�c�b
��PQ�<�''y|B�������Ħ@��!&�ā�ă���4��!����L/��^�Ϩ�[#��I���~�t�k /WR�-Q_�A��2S׎k&#>K���,5�T�'�I $�
 �R�2<(Z��e(d�sV,#���T���_���������H޸�5?3�I}���w�~�@�Шd�T�y������8�ପs�uj�N�ȑyyR�j_XP��(l #�����:90/ef�Ҙ�u�ԉ����/�S���f��!1wy�R?bǛc��kX��A���6��b�kk����a�tbï?;w�[�<
X `
�q�L�>�H��~y���h��]�6*S�@����z��A�,�'�9�ݮ�O��Ro�L�RA�f��q���
>����OUz���k�vh�:Ȳ����:"���H�( � �+%g#9��o�F�i?�����Ca�i?�Z`�O�a�Q�M4'��t�j�\M�����wй�%�H�����>����
j�_};F�I�NFҒd��d��șo)%���M��8���e�A����0��mo�ph�5ŦPeG��h33*�b���S�r��C��a��	�ܝCD�e�=*'�<xyy��W��z0$l���}8�$K��J��`��/�V��0����]���1�5a�Ѭ���A�kd�<�6�C��w���e��^S�p$Ea�*�kt�l��tS��>U�n�+T2�d���M�@6��������I�2<�I�h� {��x��{dY�)j]���)�7�tz�5=Fv����f����V�㶸Q[��f�x ��[��g�;B�B��p��ӎo���3]�@�C������g�\��*�hxܚBS�������Z1|6L�����Xع��h.$04=��֦���¸�!s[�9 �^�?qReE��:��1D�aka+*���r�Q�_��������ӷQ�ڌQWvI���r�ĉZ^d97���f8��Я�~��D��s:{�j9�I'�"���OW�lU<�w[� x{��I
��&�����X�p�Y��U?*M	M����q�v �E�s��� *�� ?	'A���a�nVu'Y(_Yqo�# �˜������W���4B�����ooG[|~����n՝��J����f�x:2�'^�l}o<�Ey�f�3����k�v��7�3?ȨR֭Ux�]���y����i�w,�MP�4�i���`:/H����EOf�)��9�	Ig!����ފCK��-=D�L���	��N����vB%+���d�l{�����G�J&�Y��DJ����`�)��o%�'	iP일�k���c����'��[ܻ> �W��?��^4�HE�3�rCn���S����D,�lʊL\/�p��.�b�&�Ӥϵ.�%�����ek��c�F�	�]īr5�wR�������R�p�Z����)�
�]�b�žYn��9$!`m?{�b�D���g0	���Sȣ�k�{��w◸q���=��t��M!���L#<5-��� q�y"a��v�@���MY&��f�ԗ��i����m૜h7��6]Հ���Ś
a?�*`�w�٘#�r�Ȱ���>J�5���h�Z7,�+bPj�B���i�\��B����f�E�C���W�Y8��ł�6��nPPŲ;]2g�����p��r�����'�.2�����@�~<l�˸1��p�,B�:<&�,=��LkNE���mM�Ӹ��^���� �A��4��#ht�pLO^$�D!��[�ʹ�ۻɹ6�&�2vq�~�h-t-��O����r]�JM D�Vf���(L�us��Ak2V��S�o�CfS�6��fL2����UZ��-��o��0��GTXt�n��f%B��������8RK\�P��<�Cf�a��X`6C�gw|�eH�݃����@3`�n��&�^I�h�-��/`�e���3t&e�(���7�@��/���f�եN ������*O	2�K�J$@��,	��]�#�M���*���%H��@Kɩ)�=,\�lGI1���Q���̟;#���#!Tߝ�s��+��RmG��+I�u������F�D��I�}���{�d�w
ʅ�����2S�'�X�a��M=�5�M׳�j�t���ھ��hD%:�Fy$qt�v	�_���֛YO�Cv��k�k]YH۰��A��ÞC�>bB,F���$�R&�Cq~%����?�,��a�Cp�ۤj��(��z_�������>�6�2����(�uU���k.��Ǹɰ�_��2Sg���i��؂�Y��ϻ3�W)6n��!�i�!۩eD��q��R F�Hc����h�Ɗ�3�o������x!�VӨm�OK�;8_w>���.��i9W����HZ8��%=5Hà�w�XQڇ���&6�
g�]�`�M!D`a�$��Np6C&�^� �x���q�~e��'���G�=�<��}��s'οW�X|&ƬU�����z����ޫGЭ�@5�g	>�$��l~�[4�v�o����� s�~�,st�>��1,i��|z��.����K�C�C�_��#��>�,��x� =�TG&���^7�M�U�⵵��j�������ZF����l�Es�
�>9>W!juY76J��	� �4�a^9�]��D,�,��C��:��r�k`A�ɰ�nT�=���Vl9�n��tz�tD�i�p��d���=^sr^A�9ߐ�&Na�N�cD��ܴf����'@Rdu˪�[t���ഩ��?/w������_����C�'y������$����Hb��Т�leC
�'.��z�wu���[�9�u�WANׅ���L�N���b���{���4���nÚZ+
ڛ�n����|7·<�ޛ 2&'�;w�ʜ�o�x'|Z{�k�#h��$��$�뛬2�H{�p�U5���u$�C8���<�.�ڣ���y��\r��
?%�e����s1�ٱ�>�7a�\1�3��f�5(���|�?.=�}w�a.H�Q3ef<��j�/e�X�u�����=d� �t^�����ɡ���h_+o����2畈zxP��	S�v�8���əcЁ��y�e֞U{Z�ip�(0�3J�[k��Ţ=� {��;N�Z��{���5��9����=H�aą��أ�����(�[&h+��PbΕS�����.����<�@�q��F-��T��׍yf��F�/�:�?�9�.�#:���_�(-�9���8z�9�A@t�q�Yq�=�!
fl\����Eׄ�d)��B�7�����FX��*t��Q�8ǒ/���y<jvK�F6i��������^,:E��J�o������� n�=�.Q���G[��Zu5�K��������I�l�8_�8)�d�A�^�G�]ҵ9�T�k	`,#���ڴJ̊ X'��sI�%x��>�&�s����;e�>bD���lZ�_z��[�����%���6�8�� -��>��@��ci���EfVv����~xm�T�K�����S$f��SoT��Z��p|�����3`�_�ᨳ��b͊������.�U�u�4��u �&vܛ�*�zH2��dU�U@�7G�L���#�l�7���O)���8�b#$�]4yی�HN��s��dT�П4�����D'��`.ۺE��N�{qW��[�w�u�cl�����������+f6L���G6��;�����B~�zg)K��f]��H�!տ �� PvKH/盳��rz���R�������8)EZ��0�a��O�G��T)�W��h�pօ^���˪��cOdP�ǩ���kpO�'�*7ð�=�
z��U 1�h�ֳELn�w�I�Nf^�=z �oBDg	2�_��Y����
K�����YPkO'+�Z���ō΅����sY������ma��/�d�g��F�~�ő'G*)?�>���z�N�Hpɜg`�+�q�}�����섟�,hિ<\��d��\ќ5IP`#C�ti*��c�ԴW�w#�z�Ћ�w�QZ�	j���Ț�ٮ��	�<�}A��`��^g�܈��S�w�um.>�o�V�l��|�b^23��}A���}�&gh�o宯3��	;�t}��"�m�ʰ�i��$��Z�-���B��M�L���%8���U�JS��Ha�7�%��袻q�c���bq~��t �Yr�G�æ �oS�H��f����hH�n{n�Qh����>[Puը�)%�2~¬�{��p�/Im4�5�^0�WnA�3Ӿ�ѝ�ubNk�_�gj����ln-@���:�uFv�c܍��*n��a'H��0�T?J���I�!3!i_
�v��g ��c��!������8�.��~��!�x�G�R��k�I.*��a�u��*fb��F�MAj޲*�3�!wS��:P
��{��2�iz��4̔_>&;bZ;'#Cin�`YA}�k�4����->� ,��U,�4�YAW }�N��]��N��Ɉ��e�l�DL�N�δ���woH�{f��O~%�
�c1��WOP�]L���Ne�Ɩ��[�;+�>\�C�f�W�@�5SnZ&C�?\Ls��'΃����ʦ�e :�@ �Gy]��PK��e�A�����[�s�W/ߊ;���rߖF�[��%�T�T�5��-t7𞫜6��s���i��D�\i�x�s���?��^�!ۏ=��cw�v��Z�v�ޤ�!f�昫��	����S�3J��}{������dY���-� F���	��(�KV��_ff�@��f���
�d�ĉ�WA \�Y���C���ڵ�W\_�l�1=l��<���_b9���V�!���*֬��t�6���<���SKl�A�/�A��ev����Ktv���QT�_�t�L�$�/T���y����&
馮�_�s�'��	�)�.:����=y��w]5p��([���#��Y�oj��BC��} ;������W'�հn��YI=��hR��*ZT[�j���,{��z�.��F/ &;�ɂe8
�����q���U�UG��5�I�܌Dn��,�����*ϵ/J.`>X�«̫j�5R�J�*u�2Ax	<�����M��}ݐT�=��G:�`�v�m���l\%Wڡ:��8+�ܦ�c�Ͽ�|�$�-�I�����W�l���o��cRs_�6��Q�V*����գ��3|`���%�֖���yi(�Q�`{LJ��y	_�?~`�@n����v�Z��[4gT(�`[��I�gk���
��Hb���i��wj���;�w^��a��a/f1ff�/bj-���&�;�3�R��eDC*�d5m�B� ˞�A��	]����{~��B���k]~�Td4�:P����%����7d���6��WX�Fd#���?i�:402i�w3I4r���@�B�N�L� 'ψ��i
�^o��NqB��I����l�"N-}-�Es��{��:^`�ˁtg|J��J����`�%�<}Ed;�f*�˺������X%�3�.l�e	�EL�ʏ7�"Y`m��֤R�� u(u7|��w����꒶��~MA�<���v-�7	t���%��I���DNx W��#*E���F�-�t�d�Pu@�'�;
$U�Z �ȷ�F��ȷfJ�LD��zKLzW.H(����w}t� ~���v�%�|5�KAϮ��_{���ͫl��͢U��Ǿ�ႇxҸ)�'��jZs���ڄ�ƪfٮ�1�I��C >>/��#�l��z>ڀ�EEi�MD���� 
����d�ī����j��i���a�Qz�<s��&Z��E�v���iNp��nP���rZ�d�`.���u�����[�0x3p�.I�Q��F�愰<ٍṶ�K�b�ث/�As�my.��9Bm�t��N���L���,Ʌm3�7�2�n����*؞�fIz���oV8Uwmc��e��l������{����`���BZ��LK��f�+�c�����H��88.w�����U�{Mn��;k3��O���)'#�K^R����<���W�)F7hb z�����]	hm���
��2�9I!SCf��e'I%Z�\ܰʮy.��F�f��Tq��׬�f�O������$�yV��aM�v��L�A��t����CB�|!M
�uK�ꆘ^�ɬ�)��Yu�L���!m��+�A�I�pږa9���e��.�K�.[Dk�,.�~p��9t��rAO܌�}�~Ɲ rM�!፾m�n�,�k�f���FuX��lƮ�����0)93�햙��ʙ�H�tW�� ϬD��E����'��f�8��%������T�Ю�4�U�-�FF cT�.���ϓ`w�͉��J��҂���[nY>֦J.��7��R�P��=z������]�.q���^��� tQ�9��Q�ig{[�w��~�Vǟԏ3k��D��W��&dITp�?}	�N�!,Z��tѯY�U4�In�P��	P4F�B�'͋=�� ���d����M���H�w��3��ב� �=�{��pC�����T��[)"�'�~@7w����%����N��?�	fH`��;����an&T�Jxq�̡�&C��JM���C��H��d{>��<�Ó���E;ե���Fƺ��)Z		܉0V_� E,�	|N:��#��qH�v�yO�����N���}�'�m����ȍ��-�Z���Z���Q˸&\�ڙr�yPK�Μ�w�ʣ6����jh_��(�'*�V&�a+�s����;��r��g��:5���g���Hпu��@�g��ĺo.�[|�Uxn��u<��~"�aOBq�� �������R;$~�����U��$�T�7�Ǒ6�$1��!VS�qQ��C��S){��D�s�^�����]Ϙ}V/z2Wa@/�C6�q�O�"�F� Au��wV5���q���<����ߌ��i�1)6S��,d��Ͳ�F��*��� �~RoBXH�M����G�{~c��Bܷ�H+��������&�z%��h\��]U�G��03�IL�y��hS'L�/��wHg�������}�w#E�6��Tʴ_�o�a�2�4K�r��mk)O�uK�/��7w��j���Z��*g�'9�Lߺْ{�}V�Qt��������}�xa�J�F��F�%tC�c���y�R���A�M�z�Ni�V(� ��eM�)��X߇;��
��2wSĈ�U������y���c�f؈e�b�P Œ�0�d� �´l�	����R~�=��7h�jo�M{� ��.%&q�8�Y?0��w�Nz�G���� z����*͊Q��2��Z���G]��Ry���>�g ����AOY���q��pWs�c�]�"�Cwg,���2��u<JvB��U���ߍ�-[a֪�q��ͥ��T��ǃ�.�t�7&��}��fO�E|3$��~)%�%0.���lIf�!hy��c�[CRp`4�%�u���LNn�=!}��.�n+E�t�-A���z�%^���X�=��}��;��S8�Z�~��������n�b+0lw�ꉪ����C%����z�	!;�e��Ñ��R��G�/x8���D�z;�9S�3���������"�?^v6�HQ��*�/�Fz`�9��8��t.BX�����έ*��1��ՂP׼o�C����dR�Mu��09cx���(��yEu��hꘚm�H����R��#�?���U2{q�.����.�Ic,A�:M�DX�V��&�<Q�e��-�h�7L?IB�C������$}	��h�V�ly V��Z?�������|6����V�U�&w^�x-XS�<w9;(�s%tW\�u�\8Zu�� X�-�k��.�2����A�l�(n��ߺ����NI��)��u
�xo^��i�iia������T	R`%��&�d�������4?�9@�x"��:(˴E|�p����uDd�5V�ٙ\���X����N1x�VƋ�CJ�Ō���0Qz��Է����ڟ	u��c���U`���׉�}D4s� �@�LwV-���K� n��`
<}���<g
��v.��"�~U5�5��b���f�"9�Hp�*'��x���1*���Q.VEÈ+�|?+�� i l}�����&Bk�V�?!��>�*@��R��r�L\�g��өT�@�H9��V\���{�O�px_ݶZ�:W^Mg�wux���"(
N�-�����|�1���͘��݁>��"�ڝ9�N��Q�-�v�8�/eq���-�`�����y|}4d�"kS�Χ~�x|1��>����x� ,��:F����Y&F�Ɖyx]���Ĳ!�O�Qe���T�׹��d	"�t3ݲ��=�b���i���y �<v/�`P�d��3�s�H���޽r�JZ�`Ux\�9@T:��̶Y!�?ċ�l-��,����ڍ9�W*�����E���L��l����KŁ�����n'����k��8�t8��ߕ8$ol�G�� T�;D�MO�<��6	�b�j(o ਅ�>0O���q5HO��U&��+�Viw�ZQW�lV'j�c^ظ�|�N�[�V�CWZ`7\�ҽ�`yl)U;M�5���7���	S�ޒ���^Zw�b���9�:'�?;�Jl�db$��D�.�A���|��P�Y�ʎ������+��R�V�@�1h ��Tr��b˝��f��em�[:#"�����1O��<zv�"���A�2��٥�>X./�ä���_�V�Y����]�Y^8Pbq+V�b�
X�S �+��q�K�A:���^�܆��&�ȟj��S_�.%�`�Ғm�+�DM��s&A���K�	��I�x�:����Lm��\����&}I]g8@���>՟����v_7<�ϓ�k@�+�}��8Z��\".��z�uem%����$lo�>A�Qt����֘��cmLp�V\��i^!q�-�\�(����g<�ذ�����Y�v`��,�_1���%�s�y�8���9��ꩦ�D��V�U�2(=O�F��G	��
�o�Ɔ��rEU�k76F6^In�u��cQ�@��,�,N*�W�*{NEvβ��)Zƈ΅)a�uF	{	�a�,�fO
���r�C�Đ�9�H�+	mMf��h"����N�%+��'}⍤�����L��8�y�|uHj½�����HC7��A�_V�6��虦>�{�@�w��e�6)���%p���4�xe����"}4
��p��(+�}F!Wڌ�D����tf3�@�z����~��)Z	�w
0XL_��pTOU_�)�!� IKfi+�J0�Y�Uߑ9OFl�ܹ-ΰA]��?�]�D�0�3W3S�G43Q�E��9$�l��
���󫢎>430��#�F���P��6FtF��Z��-�݀��e����:1����p�	G�������� 	i��WAD��:Ƈ�|�
%� �-5�L�X!Ϊ�.;�*��<J =hKwFN�|��]�
L���U�N��XV�����p� �.�<FM�i��,���D���d,����t*�K$1���h�7��詔�j�,�(�������� ���-*�!Y}D����9u�,��&������&�*Pns1���`id�0��Դ��>���`xKR�>�j����UH�U0�f�$�5U�O�R���Q��~�5�t,�g��_�N�5~�&}Ӹ�ŊHe����z�,�(��لVㅟ�e��_����}fhܟG:�'�1X'R�8���O�c߼3�sjW����B>�GH�1�vU.�S�J�r�?&q,M�W���:��lMFj#r����أT�m����W#�Z\dAJz5��_1���#f#'�����+~b3I�8��s�V��B��n�*4M5RV������J?���;�<�Q�b��.���%skz�d��ز�ĴF���̑�;6+�!W螠f��Zy�7��̭��I��ٵ�|�hs�H
�_�s*��wZ	��֢r��떈�r>0i���򣻦!�c~:=����ʈ����K F^����&z'�#_x�m�%�	��(��5|�%u%�������U�搉I>ɮ��*����;�*Gr��6���l�QK�	�?��a�@P���P�/��ۋ�����F�#Ez�5�u��8��������2�܎�ן����]�O����-z2��s �>�rW��9]L� ��`Z�w�#|Y�S)���qi�E��~��]�OJ1�C�V��EmH ��ANX ��p��>e��y�~	o���XoS3��[_�)�/6�:}������oK�*?�]�@���N�w�S�gv'��.�~uN�7���L�*���_�C͝��ŉ� ��"��<��v+�t�U�H�y��-��D���.��Q�w?cȼ5bY^�%�E菾��`^��׎�oyY���݃��.���>�8NL��T� N�Uw���edx���k4Mw֟��u��5=g�7�6)�B��3�1�0��h4?i�8�n@�a��/�3����n��wh�I8˗EkD��3��/�� ���� ��_B�(ƣ����!�5�G�+����Mo�~�w	���9��
����̉�N-��$���s��Fdm?����������;}J����Qɹ?�i�05�C�ʌ���u�𭼁�>���1L���#k�2��c�V�a��M驙s��˛���P�����������2}��	=*\�a}A��i|�k4�Ǭ!�S����M|�-Ͳj�O���U#����9���\\d�+�;�:�E}�c�����R��ݼX����xsH�8�����AS�����OFS�5_��![�'�$��Sd��� 1?$2H�:�ĳ[-s�f#�$�t�i�J��F��w"X&
@^/���c�9��Ma�ahڜ�`_�V[Z��3Ә��TE"ah>+e02ݓF1e�3�@�"ZW݇���뿢&�f5��f�B$�+���0
Az."N��\B�I�A��YmZD������Sچ�����D�涭�q�-��6���-Q,�����>R�+�J�U�Cq�-[S��Ԕ���ȗ����Q��)�u� Gqۮ؇x��g�����e*��^s�X�N�ln*�^�3~��S5i�"�4X������#�Vm��l$#�}�hh(�d����N�a�l�1��.ܞE/p�ߑ\�%X3/�m��DQo�Hb�Zhz���XN��Pwׁ��[�%B�a����|f�B�8����+��,==O?������Z}7_B)Rw��:���9&�;_on�z��c]%�h�um͞h{C�J
�5�o��뇐$�MJ1�e9i�Rd�k:{Б�^�����q� �4G�(A=rv����8���7<֎�=-k�8�!Y�nd�f�/���|`Ə�����.�)�.��~,��&��@������h
�uUZ#�q���ʱr��Cv6vA�,w�u��B��[ x���<dQU�i�Q��l$?�E�ؑ�3�C�6���ke��_�	
)T�� ��fAI�z
 ��FR�P:,a��s�;��Kt�ysl�^ �ɤm�om��?����9F�|ʈ �������ww���銅�|��J���b"�wʈ�q�1���hC.ꈂmb�kC5�I4�C��|ą�
sI��Ƚ�Dl,�齞�o4f5���gX��Z��'D��s����������+o��)�c�����]۶sO��I�.����{�hQ�V-��+�c��[N��z2����M�i~��
`�����h8\;3�X��N�[#���	���lЏ�y���+IC^�I�v�H�d�GZ`���ڸ�k���xxSK\Ӄ�Mqb,�-��?&I���.N�g��o#��:!Cϓ�Tپ<���y�'R���V�򭞍v9j���Y��33�ZHm���Z][��FW�Va�XS~��Uo�&�\*P+qy0xWyK+���/�pJ�`_�\����+��݅��=��r��}�m:i�����|�@e��t�YW$�)@-%8�2h���ּ��q�ci:j1���%�B�_��N+�?O����47|�bm����.�/��c���+`�5�q��i��1Sɛ�l�<n2�
ـ.���-���tXJ�4�VFg�yYg��Ai*
:R�?;<B��.��|/�hf����G�H��(�I�I�G[����@÷��'L{�f�c8'�BbB�&sH)�G�/��Wa?g8��g��k�a�lF�}�J�N\7�Fz��%эRht��廹�>�>P�t'~_�g��b��fNl�ag��*#تm�ۿt���/t!-I}�|�^��塁����P>��5Î ;wU`.n�˨�m!����i��ƍV�Ky���ʸ���Bz	�M�?�����2AM����S��	��=|�uo\h+�xd�r��Y�=�K���n�����GS��k.�́S�O$��ܜv��˷���ď0Xr�ݠ`1�M�"�=zb!e�گQ�	�bS�߲?�ڟ��OR9����X�b6|3N����ŏ�����>�ם�f����~�-8�A�k��	.1��ԦC�ma���c,x�ݎ$��L��}.Wzl�PS��@[�15ǔ���V�z�b�G��:��.��K�-�S�P�ۊy������z؝��}�F[�L)X�P"��3�jb�Sq�����;��t��q,v	3��ڱfOS�S��`;�3�A,�⸐��q��8�UUR�m�#t����E��(������ �h ��4L'�kV$]��q	�}��0Ss�!�����3�aԙ��_���xBKf�㒩�P��LC�-����]x��,Њ�_.��YW`�����8���)���/�����R�^8��AjS�r*9������ޱw������V�i�]R���V� EQ����$�^��EWs����;���1G9��������0�7Ȭ~�c�� v�c��n��R��V��ڸ����6�c���-t�e�?�C��L���oMT�Ձ$uC��-s���&ݥ������V��Z9N��iO����@\���F9q� ���.K�e��|{��F7�m6�BCŧ�V�>�����e�&̎�09�`?�f�N,TȽP�:�����h;��mte\/a�g-Fߤ�c�~���e���OMu���� ׯB;]�c���W�r+?c�i��`0�u��GD�J����m���p���Jo���x�4����~�����SK�
J��j�X�|���3ڹ*�@�&E`S�/S����z+��Ub�]?R���4`k����r�T�UY��Cě�<��|���"x�5����K9�iG�	����Df��.Ӈ��9�>�
�KF�G���gl�\:@�%i�e'�cmx�
�5[19 �욿+-i��]��P����@vie֮��b4P�J�s���<='�nh�_����/����mȃ6�r��@HJ2��lP)E[/ �{'��`"�Zoy�i�`q��	m���d;�|�(��0P�03N�E������M�֫1������^f�|�b}��TFρ��	����3���������[XF���Fؒ6��O��/�ӽmߘ+m�H�\��t�; �F���&�U�X���@����2�rRx�v�
���8��WR����{M��ה����7�}���8*�H?D[_�9���v���.J#mY�Ϟ7YlC�lES,�q�吗 �"��A.���F-�l�yc#U`�b����3�сƮ�!K�6}H[t%�l�|R�l
���n@�����������i�D[��^ (���ܘ	yMڈ	M�O�o�S6i������7ʐ�e��re�ΐ�9)�?_L`GB�jVr�0�#(��Q�w4�� p����+�|�������>8�5W��%#��E�O7��8�B���R1�g�Ӎ.�ș�oy��(̍�����먄��dƞTm��@OƄ6A��5UM(R��C��rwN/C[��˚0��}�m/)j(�Q��F��\�Ą�B��B���dj-���*�pOY?���J���#�0��Rq�j�b�6e��._�X﵏[��[�����*�wu5ڣ\B��L��;��g�� J���_4��{Z��u�]CIt,�r����?�DR4	���i��
���ִ��ܗ���(�-���Dq&H�����E=b��Z�7�����ζ���"es���x0��BM,��q�4ݴ�O=1_�;qezS�&;�X�Vf7C��f�*�`1}h�/;	/�i��2�F�_����q��a�1�'���4�VV���Ax�Õ(ׇi�PXD���;�'�J�πX��X���Ŧ�yl���,Tj>�*c�M�p�x�d�Q��̐��xc|V�o��Vf��^[Ce_MYw�F�F�j����!X" 0�T��g3��z9��bE����a�y�q�e�^^P��l���+�$3�R\��h|:�\w�7�Z�R@���)LL'�>t�e�A]����ST|�mG��fDX�[�x�ŕ�g���_�ٙ���u�q����3��M��W�@B���:g͖`Z���O��-9��&?Z㧴�>k���D�y.^s�y,��ד�b�gp�y��)�������3�} ��q��;�h#��k]/ቫ ;m�KZ,w��8Q)�)��	�q*%��J�X��V���L��So.�iL	`��3*��;Ԃ���O��؂�j��Y�&j<�+�Q��|�X��R����Oފ��P8�,��1f﹀ܫIi�Z��&b��>SL�>��¥�?��\1%t��;��.iE 9�lZCc�F����4���QpoW��ůV[���*O��6�7�%��*�w6���"�%F���̘>�{$_z�Ӂ��+�6A������=A���C�@������?r���~W*i=�(��+�1p���Õ��_�O]���!���P��@�A�԰t��(=S�f�=�#�Kհl��&}� 
�kNwZ<o�m�9�OU����hr9�����\E�B�>�����Y3T1~z8M�#&�׫�K�xAWx����~�l��Wi �l^a��v2��7U+i��
yNH�R t��u�q 5����R�ȖPu�2|Ux�t�j�M|[[7�-��@�z���O����j��F3�o�Ɔofr��<��+7��-�<�p���NnfV�h��K*����+Uv?��z:�X�<��f���$�+�IezᎧ���`:B?x��3��G?_�DvD)N�I?�ա<@�R߯�2��4sD� 1����",�C���*f��-I(�I�l���������v.'��
���Oo|�^G�NA�Q��,�ܲ5!�s5���<p'��0��	w
W��bf��g ����U�䠓7���NlD� �yH���=W� ⏷���OVhnu�K��i�e�δ�/�rM!,�X����M4��)���'�5=p�+7	S�P�^���n�0�ޥ�L��	���3ba�h�����T�:%y�g.���P����Z:���<C��x[� �f̛��A��H�6�"Qq��ҫx$��HW6a��Lhϕ�ޚ��a�ݦa#*@�"��}f�9�X��	�g*� e�o�B�=�`��ah��`f0j�qU\��z�hn�>S���ˏ&{��� �c]z��Y�M����v�C�$��0V��@��H��#B����0�Q�>�����Hy�S(^�&�E���@T�h����DI�l��2�Z�"6�8a]�u7�V�u?ҷ�e:!O¹�~�7�X�L��2KCe�J�m��ێX��a�+[�}O�d����<Ί������μ/��IXm1�[�g�s�[�b����$���z�P�	�G|���'�Hۀݡ�%|��I��ȱ�m��TO�������L�XhAǑM��U�fOSXC��i��ds3��G�S��H�r���s��E��������`@�;��Kv��S���:'ܓQ]d�����2كsN��
��MA��°�
1�w�|�[sA�~a��H��pP��esW�V��<�
̕|��%�$��8u4���pg@���z3ۅ}�X�_�z���D�_
�Oar*�w��VB��Dk�A������X�"���;~��z�"Rb
��!X)�L�� ��*;2�35?��n����A��wr��������ۼ�'"W��ϱ���\=l`�~�^SYbGum��ZG���o�6�U<��k��瑸������jbOf?��sy#�X��ǶmZ=F�4�7#��h��QRcӣ�/[��` ~�s���5,�"#Jڈ�yuaO��3O
����Y|ن���W�M��o�ͬ�\��)�����G-�.�=�q�^N�9]S�b��9�Q��\N�z���a����E�{+�>e�h�oW;��!W|�s1oR�tr�M�YG����s�L�i<����Y�-���Y�=��)׻�Hy����%�79(�	�"V!��B���F�i���x��5��-7�|L�������Xo��B�3���/����EbT� 5��/��5{�Ztɣ8���'wr�-ҷ�!q=h��ȷr�D�l�֣�}7��|j�����!hB o^@�4��baOYR� �0c����_�M�C�j"̀V(���`K���ۼ{r���|'kK�������Y��_�tT��W��ߣ�� �0	������
����U����>��.xH�[��*vw�r�"[��h7���nG;ї�����$���4�z�̿3φ�ދ�l<x�{��,����E�[ՃKŔ��me�V� 8jH9C �{����(G�Y[�m���*M�|���KJ`/�ͭ�p���zN���9�����Qn+
��Pa��y�\�͋��ɉ�������"�b��k]�s��jo�Fe^%]3-jD�A�V��ڐ�NgT��w�|XPD9��.�#��*����`ȕ>��zl�YN���d�����_�)i�A���l{2�ʆׂԼe8��pT@�׷�����T�-|;m|:�3i��z�gSV��57�o�1�B��^&�w_�ǳ�y;R��I
d�6x~"Gٰ�ZY�#��@�n�e��#�M���)p�P�f3��Y��h)�K���ƹ���3�7MͤA��&���o?j.�	��ՈN�)�������ճ� ۩�V��WT��M.�'�A��cL�~fz�(�6�-$L��3�'���r�NCU^�	�ך��������:~�І3��UI�`��p������A���B"�H<h�
�+�B�Gu�T�V To��7V`�̢��,A���z�'qٜ�w,�=�Z���:�n�%-*�����I�g=`a[8�����?�Op�0��4������C�FO��h��ɇ8FX�<���UƎ�؉��������r*<b�؛\7$
�م��4�kb[�Jq��"]��Y��

�c�J�T��)�s�0Mޥ��[�=�3!w�ó��2�1�	�a�WR�ࡁ���Ǳ��.���\M�OWM�<�=� r69�%ז�c�(�r.�(wb-Mhw�N��"�a�w�w���
(�~@Y@�Ս˫���(��!{��+�V���7�,aɋGvv��EĤ��K2Y���,���k�>��P���Hx��6���Z���[uo���o|��������y�w���Bea~��2���2��{f(}~�t��z�0�_ꋒ��1'_�P�yU�#�`�<6�Ȅ(M��,���=�P0ey������	�WK�@)�K��ч���$ Ǩ�Ae���/d�)d�9 ��PQ�}�������G�����4e�p8��@��zada�;vp�=�sp �خ#�dv�V9#,�T�
dk�?��瀧៝|ek�Q�Gd�R7�]��xY��Q�ȡ�\�Lhs����[���(�g�W�p�7���~�6�nTz��N3�|������H��8������*T�hʛ�M?3�74ٴBH�c%�rs���V�2��n�XYyX/BRe��_�WE�)�Ol�>%5��<`��PFv�=�~+�s\ʜ�ώ��R��9�sIy~:��N9������i�y���op!��DZqF�I0y\�a6vor�m� �RP���e�!�'A.Y�ᦇ�ן���ib�^�I�9��7�#fyy�yP��S�ψￌ:)���rЙs��|�"��BX��s�ٸW6�:|3��H+kQ-���9W�����7���@�f���vf	���e$ �0���}#;���i��8��'������g4
��k7���?����stw��ڧ@���fIV�D��<����Z`��o�vKM���eB���������R�M�`mxe� �e+�%�k�7�oL�.лo��~�A�E�`�"���i�URq�u:�.n��9ĕ�u�	&����5���ĥ!�[Qn�x)������͓�pz?�FO�~�i�W�E�R��#��ZPz6ɨ�é��.��ڷ`��о�SҜ D��9�c�I��[��)����	nq7ƔDs�f��e.LY�!�DC�m=l��m����ݫW��dq|��A������2:R���;��O	7�e�_�V�,uYs�������?���5^�Jv7|�� �����՚8�?.�NZ�T߀i��{�QVԍ�V���spc�fz�P��M�H3UHX.q�U
�n���������o��~H���h���`��|�׻ ����r��ᤎn\�g�t�Ψ�B���}�+ģ{P@�1��@@N ��ck�_�um�q�:�����&C=��S��2��M	V�ˌ�'f�p�wŢU�]Q���$��&W�ݵ)�7�dp2�^L`1�3.�H��69�C�
�kX`�ZgR2	�%H/����&�yBD�	��B\/7O7^R���@���I�x�1��옠�i�Dmˌ�� v�Vi��10u�:A�7�J�z�UX�.�t��ֿ7�D �
�6������W4@<MR����1Af���W9˯��)�9�>!�z��듿8����|0�ӏc<�s�
ؗ���� ����t��&3'��d�,$��OücsT��p(��g�0��*s����	�^��+�ۣv�}�k�j$5MĒH���!��_�u���<'�@���ߘi���:�����q*	����S��щ�9;�=�!:�����8�V�����eUT�BH��0���p��+��*;���FI���MS�啂r��l�0��_��*�t�)l�o�]��|&���w�.�<�.�:8��*�&a�X��u��,E~��l{mm���+��qi1N��,`��3��:���i3!���M�b�>xg�)z6� um#�����"�>й�(�{	�2��� �3"wTh�\*�#	���H��U��AG9��4��Έ�7܌kʝ�ta\�&���y�[0��,�A�yĈR<��^��X�}u�
 _�<m��sz�@�`�~��)�;�3�&~S�AFL�a5��hk���fs�%���~�<O����ہ���A:���18����C�wJ�����/�6/�W��5L�n�XA�=o�	�6.��������̢���	����h߱p������9fNH:-�e�m��B;zH��"
�P ��"n�h8�74<���}O���1�h��#K���&�� fp)$u��\��i�����o�1��}�uދ��m����$���t�R�l�k׍m�}�J��l�Q�"5t4��X ��`�;�_���
�K�%D
�Чc07h���T�t�6��k^�ms%�����ܦ�>�Cw�8iF��i�b0]��<�� G9/�+3�'�����]�efڶ�����o�U���!�'?$�7A1���?�fȱ��������T��k�L���8�<@D�+:8���7��OJ��_j=ʇ��N}E|��E����
Tp\l\�ަ`�K*�����.T��R�����_]��v��7�gsX0Ku�|�Ԁ�u�F�b��G腅���:q]��N���(=�oW嫜��q�m�>䟞������Q�|����yƮ)�@)�^���_S�+��I�Z"TxI�����" +���Һ�Ƣ�6U<h�xx'��w;���p�%��QHC�E:��ҏ`� �O�BP7I_G�����o�;�Q!}��&�y�E�x
�h�2	#ٗ�浌��hO�<���;x��[�i	�[�e$��u��\9�� �E�b���־Qۍş<�T��/R(=��;홙�X��	�K�l���eRG2�z0X6��W��O��n��$��_� ���F��O&��f31F��
�܅Jy���L���Q���t��rY�n��e�n��O���6Xm� ��#-��K�����]���à��KJ�k��#qI���8΢��;�ʤ�X)��B"�p��G��q���	����RW��,��jKL�I�6�*�Q�J�x�l�xR��U$��Fi����7�-�p���G'��ȧ>�LXɝ��~%!hq	f�U�K'-꧆,Qzgo�b>���"	���ņ�s�"%�P���9d`��
	=|?4���QW�P<���=�v���٢p���"z���:�$�o�ET5H�ݠ�����N*&��F�&���=��EE�����Ae ;��V��R2h�VN�
+˷��'7��hB�I�ì����A�`�@�f��{���~ ߦ��G�o�!j�P|��63�}�.E΍%�Wxb[�)���
�r�A�x���\�B�-53i�Xڴ�R����SU�>����uG�|��#��az�~a3�[Z/�7d�/_�}�v_��(�W�<>FD�G�p���oOz��eP��c�"nSky������<�s"�����T��[\6����X�G�� j"oR����f!7VM9 p�6�w���oyR�a�p�,`KbF*��6J��V��6s~�g"��.ء��K��Qk�.��aǼ�7��w���<Ox'[�*�2�[�6��hd��wK$�V�.���d�3�
��V�T|��
�n���Cp(�~�$v�缮���G�ҡAYۭ�4�y�k�62��#��=��7|��=�9�u}F.N!����p��[o���o`��y<K����8��g6/�(���Pd������ݶw&�zE2u����*�����1qv@� ���,y���P�,{O �)��Фp>�5�>�������/i�KYY`�N}m:.���A�h�i�̪_����G�<cQɜ����ԗ{�[�Lo1���W�'�kwO~�Ŀ2�7�(\�L۬���VĢ��7v}�:�;؋0I��L�G=�,��^g�L�s�#��5(+�Ǳ �D)���q. 6��f�^�؛y��ǁ�3M�.�'U5jh����*=��0��t��X�*�b�,�/�F�@Qc%� UD}��r�;��G��!��(ı?����q#�5G[hX�����l� ��������u�Ш?�u�&�+�O�7�hsg���eq�a�L"y��:�Nw�D�i{׎\ 
�ɹN<�����t0��OQ�� �A;y��)���ZyOd��?LeN��I��벖��1y_)η��/���>��4�1�����5�o�XM66�P�e<��ļ�U����E�H��$58lV�|X�ڴ��S/ �F����_�g %��D��jo���.�8MA��e�\2|U�sϷ��Xz�hZ*����v��K&mB�3q Z)��Q����F����N4�K�����>Z�4x�J���:���~�Z��.�c��sB�D=p@�B!��Jz7JG�DpzAp�J�Ow��ҕ���,5�f���7����1���������Q_��������e��r�:&�i�_�1I�icS�F��������xȞ_#:�S��K��}��1��f��)�h薵�@r��ꝣ�����~��#L���tn�J��*���H!�����⚊�N0XM	��]ã��0W�r����ʎ�����@7��s���dy�A�02�=i��KO�ӆe�>B����
��ù,���p�(�!��-���s|�!�R�rm�wX5��O��C�m;����߹��g=�L��p��������x%�W~�ɿ���JB�Oc�L�1[������ү�.卋�� A�N��>��Z���S�ze��wi�/�|�K���9�0W\�\�Z �E}�6�C�]����45\����jw*Ϛ�]Ij^T�h��'�ʩ�j0�
1h��eLg �����Ai���.���4q~��O䒵F�J�!X�O?�N �Ò�K�E^`B0K�<��<&MS��O��<T�j�v%D��ฆ*�2����%-���Ů���>�a�r��_m1{v�R㧾��R����.v�yτ+�T�[~�!;�}�y�bW{�|�%�F}N}����~,=Y�o�aR���Nu���u=��PIl�4�P5�g�	�)A�U�ȃX����Z��x�/|6E� ���i��֌��z��N��4C����;���u������Hhb�HW2 1�ܧ̊G����P|M�斵��%B����m�ڛ؂8�%.�JhkRyo+�x�-�R	�,yx�V�cv� &v�*�N'��[����Z�����k+�RL6�yE
����	x�*�Uf�P�&�+�Ň+�9����cpW;�ѱ�3��J�9�V�7D|��$/ӁO�~̈�[��P�Ȱ��Ry#�����q�.��5�a���h̖�D�>�$O �3�K��"s���7�D�jŕ��DK�D!'��`ߊ��{����(�(=7=>��@��pZ
-��D��+Pp��K6L��n�v
&B�ls��-��1��|�/��D���mV�385��,Jߣ�C�����^�*Y�d!��#�Ȭ��ةDɹ}�@KDvc�E=s�9��=��;hb-AӰ;4����^�ZyI#�%��
�G�FG�4B2G�c��/\�?�?��Z]��Y�;��.�Gq����e_���ǂ�B�]c˫$����ӜhƝ�:n.u!6e �6C����}	����?��dlWA�O�H� 9����H7�.�0��������b���r�[Vm�1yR����Wr���j,�]�bm�޹���l�}F�hMpڟ��PVE@RY?��ă��s-�ק���"��	 W7C��#[y�NqjW��E��O�R��VXe���N�����O�Q}t���'*^���D�f�`=�@�R�=0x�,���U��Љt�49`5v�i_���(�
�F>��[�����d�S\�#=J �]��R��l�AK��� ��܊y�M���+��#����(�L�4j�x���_�AFEo�]�Aɲbc��c��H�+lt!�Ha��b���h�m��C��n��,��=�C^��
$<�X�^�ͳ1�8f�^[�h��`�Hjh���ԙ�*_�Ԟ#�Ȁ�Ӵ�"S�g1�=�%	{�ࠛ��" �vj�$�7������-�"����iE--d>��E5����
�o@���nB��lN�]h���DF6�[�63*ڮ5�v��%ko"����Gg�\=�G��?>:����AJ3�����RʼsG��yA���[6M�u����C�7�*)#7 ���5U���B�3K�p�&�_���l����w*g�;~i�t��kT�I=�Sګ�V�^R̴2h�+[��ѡ��Z�ϗF�!�����/xM	*�߀O�i\�@�	�����G�h��Y�M�Bm��2-!4�#{ :Pyi�=�B|�	�
�S�x3��|k�滛����
H���o�Ղ��8vH��Ƥ!�E�?�#�'P�R��'?�����h�8�7�F�ؿ57��$r,��[�v�<���{|�Q٨������yiX��B�.�i����(��'tȱ-i��i륑�I�U��ڕ=�� d# N��w�
� `f��V<�Z���U�)�
l�Bh�RC(�/�#<�iQ���qk��0Q՞ڗ���aA���6�'[P$���y���^
M��W�#����bzL��2q�����qs�aCJ�#-p�Q�1��D����5Ǆ�q����}N���.���J���; �u�qv���@F�[֖}�%�"���MaXF�xeݟxXP�Ry1��}L���!4����	~��G�VS�|z�[�U_�R�a���|L��!2Y�}�K����=���JШz	NB^^N"� 	V)�T._�D����V��p�o5ݐ��%�r�ޣOuu �:�[,�l��q�F=��Q�y*7?�뀁ξ���z}4R�_=�b�����&�٫#����L������-��S0!��k�a����}���T��.jHI╽\#�_��n��Ɣ��ɷܸw!�����m��^����A��M/�yr�k��cۈ�J���ǵ����!��Z�U�O�(�3�qj�*v���}�Si�5(�P�'�c\�R�!�k.��ߍd����P8���XoF>��L%E��o��n���M�X��tZ&��8h�y'I�th@�n\�ڦ���78�g���#��S�#'����nν3��L�i@�N4��6m`��[�I6�Q�t|3�/=mS���>հ�KF�4z!�X��ژ��勮JpM�����T�oP�ݦ����tތYukI��x��;�!<���}o��LN4��<�'<���2���Uj��L-&T�srHE�Ы�c�BZ��,'Rwf_r�{9J�K(��Y�o�V��#Z�xS,EF�2��f8ej�(iy\鄲ٵ/�t{��c�'����a����f�56��=��ƞ&D�F�+rm�'OS~�	6�D��'j�wW<u~�2�Ǩ`*�v�m�K7"��XV��5i������h-���R�퐎(���ەhZ�����
�6�9D�]Y�����ʬK�om-�y����k�8�������ecX���ѵ����_�����d�7��ٛ�@�j@t�J�|���Q}� ;EC;.�ё���R�:����Մ��zA�=�F��5ڲUI���p�@� G�`.іN��M����S�qbAv�
��N2a�@��)S#�����	X#��kłb��x���&��0�Ӄϔ���SJ'�=|�{�g�!��'@�ϲ�y8Mj��`]O����[�B�@�Ί`Ze̕��7uuɩ����y�q�0R���;�����c���I������Uw�[#B
_�.�����N��=z�GT���a��������.y�1��7Տ���� P.傖�f��^���.j�-���] �S+n�'e�<�^[�2"4��oӎã:Ҳ���5t�ѓg���3z#���ۦ��|�k��@�@�$l	�XOgT�r>��2�>����,�X�R���n˪�
��Q
�mN�l�d�6P��K�!�C�j��N��<ZM���t-U�r}'���d�9n2�XO��S��sr%�g/#�ţE;��Q� �:�I�ѷfϛ�������ۖS�	(��5�C�
�)��t��U.�ur �G��B�p	R�qͽ���%�l�ے�3N�wJ�G�5QQq�Pv`L_dJU���x�I)���g����dL#��	������e,`[�ٷ�0HO� B�wz�懘�x3����F"�2#A��>��$.��Fk@�Y��H@
���>�^�@D@����T�N����]P�`�IZb%�{�����)�;zt?����O��ٗ�q�P]F� �h�WG�Xz�g@y&H�%6E�#�G�D��gU�O��p�?����Β��R��?�rZ�R�)S涺��/��-s�}r����J�2GㆧC��@�X�#[e�����4�?;`�aɢ��ZV�_W>��7ˌ�Z�.+Ď��-�.U�E�3��������Sg��m���ޔ���Ċ�Qֈ8��Y
v:%�U����ZABݣi�

��m��cGU���GZ#��8m2�vn
��0�68�Y���M�I�M�XXJ��UdƠ"R�r@5m�k����M�����f�xA���T����� ��{d�5]b��b�i-��#��q1
\=ݟ�c[�lG-F��OP�K1�G?����M�
^ �/:-�r�/�Ě�����@\4�O�:L��/1n��3�Af�_'�e*�����%b��B�pE�(����0��������k�X�@u!��=�&z��ѷ�*;<S[i����a�B���Z�R�>� �{��"8�bA[p��Q5
��e�yt\H*2D�d>^��xl��wnm�ؔL�������IQQ@�e����.�9��%����-��U2��IT�dVϺ]�)��R.ͯ��/�4�k��fDڮ��ԕJ�b ���A��;D�������edjQ`A��(���� Lj�]�ą�r�UC�v��C�Hp�-b�$z�`�n�+h�R��Į�#%��7W����W�5��iR�όY�ï��n��'Ȱo��[��wZ4^���h�����1����SPl�+����d��8�g��hp����v��S���!wUkx����GYÓ~��)y�N��B�����1���̩�I�7FZ�c�¯M�0}!��^� �< �i��X~��؎Խ��C���<^���jC gxt���D�Ӫ��w�р�b�A�8��r;�n�����X�mHM?E���0"B1V=I�Ru5����P4�����̷�B�~��2��":8�%�5�EGxN����>��n��n��|�7z-<��TK�����9��d�7��p��:�XQ���f*��������-�~,Y�tiE����DH2~���ZU���8>ø9Nv�=>�e�嗹�'�V���h��kۇ���)�k����L��������,c�zH��vǆZ��k��A�D�����\�.]�b%��.�/�&�����Iygs$��eqiF�L�@8����#4��J�&*^��Ϩm�^m��?V���]׬U*��/,W<X �C�����V���VCXe���P�?�>p�>/娗{9S���]��6����Jg�B*9��z[�T�5��2Ӕ�*i2A5�[�vY^m� 
���N�y�6"�yKp_j@���C��-�4&%����#�����@[��߱�u�R�Ҍ�(�1��N|�K��<���k�J[�S�(Z~[!�Β�M��
\��|,e�g)��%���TX@��,Z!m�$߇Bjo&��7*qG��%8?�H7N(��C6������r}tX�'Dm�w�=\��X9J&�微�*�eW<\�%�N{8�[����7�X�>r��%���qt����
�¬7���։�M!��`��-#}yR{�w�8����E�~�V�^˼=���ŲG����.��~��!�����-��}�1���O{[�O�{�ŝ�&��|�{Ŋ'.E�CJ'�j�4%we �usҬ��M�s:8<ܘV�+]�(M��RNR�� �P� -�zFD���6�T��ժÏ:��Q (�ͱ�7��&̲�S�o\�:z G*�V�t m6eD����5�79BM�ˉo�A{M����U*7�q!0���=�䛌�V-p��z��ȑ��5��
�����qK�y�N�?aOkJ�B_�B �=& �߄��y�ͻ���q�d��k�k-��x��p|3�2>��=?��3vm��MHA�ӭ�.�!�fx�)M��4�`�����l'l��������RG��`F�B���z&Ǒ�6��v��gn�!�(H����#S]�����J����g�W�A�����u��Ǯ��d���'@���g���~��d�z:�߸���j���$�)#d��%+??
������A��3�L����D4i��٧bnl�\�������u�ڍ�ʛHi̔�;U
/����z�5�U�����X���q�&�`��&�C��E7p~V�n��JOI�:���M������V?/��a�������מ#:�>��&�� ���ד���b�N�M��[6�Vl�æN��T��i�1u�1Df� �{ �N���;��)yU9�.[{�݌�
�dBb�\���{3�ho��Saׅ�0hϴ��.?�T �<��KZ�j�Ge�����;2}��c�4���I�N���i�F���J}�9��C��G�K�P�S�l �4��iG�f��+Q"�<�F��\�3��W� �1ax�d���B�L��U�5RX��ȓ�O��m$��ft���y}���B�����O���SK��;5R'`A�T)a����&��.��5�$�X��ꖗ��'�z��M�
�8幊�������L��_�%�"�&��b����Vt'Z�ή�����,Y�0� ���"H��5P@o�O�l���-s�V�|<HyG��S�&�~�+������5�כ�;�G6~�9E3U�x2�N6���G��E�A��sRnB|�$=tmɎ�-�;���Ͷr���!\�������|�C�L�~S��Qq{FǛj��710Cہ;����0J���Mc��/+��+�h������Mc�\MG�	�T�Xs��;���Gn6L�m � Mg@��f��|�<�>WgF�X�xó��(�]�������Qyz4����t.O���3f��a4b�۔��/�Aj�d%-����58I�J�0H�G��g�롪�xG�"~�|MzE�)���gw'jzfc��\���=�\�N<�v������¥ �&ܟ
x�;���3Q�~O�0�V���9�.���?��ˢ�������k�����ks�eg���7�q>��9��$�Y�l�r�sE�]��NSF�Y�����Q[X�S�����M����,�Pi쀰���RD��f���~�����C߸l���4Dd�.fT��av@�չ�D��H�K�2�&��tS5��
yF��6��TG  ք-�}.7oPF��6
���U����X��F�w&���x����O���4�KF�3����ykq���/t-�o��Lt4�'5OشJ�/����[��@�\n�2�g��'8/hWҲ�8~݂ ^�&�f����H�L@�L���îU�ї<S�iA���Ti1ǣ��� Q���B��ƍԶ�Z��ݚ�	�N-NM�s3'��:U%=@>l���~�]-|��c�cS���_����2vrߊ>�}/�I����!�X둋N��-_�E�Q�S=�O�,z�#�(?;6��@�Vb��HR�{�#V���M��1F�K7L8�t\8��V:��!����IpN�`���YB���/ᢉr�]���p��T^]!�X �����z�>����C��*�8�5M�؋6=T:����s����r|���!r�J�����D:�[b�h����EV\Ъdy�;V�r�?��s۹ �RwխTB9n��u"��Dk*�lY�T�O��*Hs�t�jf�i��jTgL1�+͵�=)p�w�B��	%��@�P ���,��2�y8����F�I;�%��;	�v^3�K���N�s?����"��_X���g��/n0���2L_uy�w����ڱY��_������N�,�����0!	�s�n�4I�_�5+xT��80�њ*P�n�?��]g���X�8��Zw�˻����{�7a��x%n̿6Z�n6���-���6t������1�4����y�s-������=\�Qpy˺��K�) �y?�RgN$���LQ�4��z��	��q�R�U%���lNSJ���r�]8����f��`��~�m�1Fw�@�#��]j#7Y��%?�oωf��28��\-�U��E7�i���^���l��!�gu���f/kf��'&���s��5?4�9��#v�Yf��L�=^��e�|r`�
�%M���>F���}"vw}R��@�eDe�'�Y6�`\���n��pb��̡D@�8����.ć}��+��r7�zwI�`���ճ�[�oĦ�s��ją�^\.���ά���lhpp�M9+�î�XQ@�fd<I8h?�c�)��:�*��$wC����|$V�������	^i6��N�"���˓��b�`0RAÙ~\�"�hs��<�KC��t�����П|�#�(I'j�	�] �\��M��5����0��S�`��Wم{�$���*�1��`9�+��j2���SЁ��� _�c�M��_8�g*��PQ}�'��J{)'E6X�W�:�O:?��u�k#�v���_�B����mYQ�О5�z�^h���Ҙ/GS~߲}F����r��Q&�PO����`�4QE�쥰�,�1@w�gD#8�n��u�+�9�1F5�;�M�w�i)؀c�Ь�Y����_V$�(��o�\�S��� �����+� F��tk�V�nx仄�6�f;I���yj�- ѵ�uҐ�|6��x_�V�u��$�# ۞��We) ��T�Q�^�=�ټ]�Y3�����#�<��n�=Hd�� 8�4�<�'L���{r���IW߳鰪�ٚ��%7��9��,wur'���e��I�<ՁmRʷ�(8�q�+�1�G���n4���0�tw/��1���4�W��~f�z���� ΤWVo�9X��_ٱ��ʣ ���HA43/�ջ�$�e
IK~L�(��~h��Y��^��9?3�ux�{�Xb����D�PjF���+�D>L�Gh�:��L�f�K[mn���\B����H<������7�9�i@���?} �[!�dK�aG���v���J?jv�|�ʖ؎W@�7�
�b���[E"���8��V�3�܋B�� xt(m���V�x ��Ԁ<i��ƄT���kM���4
~ʅe-9�&���mD��(���� �kX@b؇��_�:�0T �\��m9�/hy��Ƙ<��"P������+QGRM
 �f]k��.�VG�X?Tuз�X�f������� ���	<� ���h����K��q¬ �.��=EG��!\�I�])����EN"����`ܦ���L����B��Gm֍����	�o�Fr� �W˅ː
Ɲ��}p��}�����V��7[�
�� �m�����d�����м�����g��^;P�&���kBf�R��&�&ѕ51����>�6�����x(������_��^]���zB�x{�`�,<$?�Z~�Cf�}�M�1W�_��-8��M�%��k@��������!}�-x�����s��n~�$$L����	�t���m���1H������$|�x�I�Х�`!�ɓ������H���q(Z�*��aL�.�A_v�P^ВN�ʰ�'iD��F�����y��}����҇��U9]�9���%͜�5��C���I�u_A9q��VZ�=����W����'�+tp
��	7�M_��$���#��
������;;���͒�Y����M:8z�=��49�������BP�s��ZMf�&�@8�����l�;�2�jeN3Ϝ�V� CGH�������W*�ޔ�O��[��,�5p�� >(
%KW$)�c=�EՀt��
�CnO`�%ދ�V��
Y\��[��M���@�0�Ƿ\�FW���>��y��P�0�;�&��JK��<�I�j�h�M��F,�3[}��p;��
���ն�+F�*���=3����-�&{���>��#����&�!ޅ�_ԓ�X����	)uԹ����5���i������y�OkG�_�hțƮ���Ǉ��x��"Ĵ�e?h�G)n��-y���$��ܜ=��G ��4]����v>��g��O�C�QՄ3���j�r�b��f�^z�xX>y�Sggb! �ә�9���;���ފ�2�� [uT��e��*@/"BK����v7i�48,���U��)ũ� `�\ΐ�6ݞ�u��?�)����4p�������p�8ҵ<Lcr�E�������Q��R�DC�#sZ��;��(5�=���k?yW�~�!l�J}3j�����k5DCz�	��ٻ���k'�BP�W�n��CE���"��q�r1��Fǽ��Imh��$�;��(�Q��U$cL{8���ao���M�Ȁ4hC%IU�m�����B���cE;�j��+L^��K�䉷-:�c������~�_%��Mٙz��iW͓ڡ¿�kwz�����׫f���2Jf���Z�sx��:I�Ǉ��X���"8�qT0�s�p���O�7L2�E�Xr�w D!x������ ��ck� �ꦠ��i6ɵe��j����f�]B���%x��D����i����"z܅n���>9��+L���$�u�|������m��\�˶��~��h(�+��_9?��KG�n	iP�e@�~AW���<���ĥF��<`z���OA�c��,U�t�z�ԣm��Zo�?K	z�8}_��s�R��Z�	NP����M%�T;�˾�N���9�B$qq�lV<�ؾ�tC��K�$�%��}^��.$,�I�R��.2W'p�q����L������BZ9�O���3��8$\<.Ld ���%�Y�-�aͿBi�Jֻ������a�K��(2d�������B9
���S�ż\���jHn�f۫�x͘J�ig�>Ϯ0]�f�"E_�S-�eiJS0������,�L�qג�-�Y���P�H^�q���!H?h�eqP�Tܔ�~���O�Qచ��fCʤ���Q-�|�I�����4� ��sX��^����2Q8*Kb�3gJ��F�J6��������%�1���WUY&S��G��W���Q'�A�Ӄ\u��5.gN�~�8|'.?x���_�h���Q�/����eM�I���?"Z7lt�����ڐ����;���f�׽���
m8 ~Ε�9 ��lQt�J�?6>����f&��<��^k�� �48����2nd���g�)���܍g�)�fp��践��x���%R�,��#�h}н�<҆Y���j+��H���u�����r~��Uh>om�~U�p�A���Ns���)�ar�΀��B�B��U�2�(]-��}�|�4o���:��O˟;�_�Ub�n��17�wEDw��3����ք�Qo�
���QKT�;�-E�)$�rX�N���z��Yz�0��o�N�W���l�N4m���S�e�YR�v$�#
��֩ �_��]�����M��ZE�����I�[�@�{��Z�E
��*ܣ"!������]2['�ل��h�ᭆJ�5؀
�kq����7t�ռ���W�PćI�5R��Pz�u@NYVw������+�޴hMv����qwf�������]N���5�b<P�ל �J0w<�~����Z��.��2�6E���u�W+R�4�!VVQF�� �en�֥�±J�R6�L�]�Z�Y��hY�h}֩�ei���w������5�_	�Q��j'�X����F��>	[@�P�YZz  ��"�d����9p��ܰ%Hq�mf�\w��|��8:i?bH2�}'�����%Z-m}�X��n-�o�/��3n��2u��6٬�D�& :����,� Y��6^I��Y�7T��f�Ez2Nd�D=_���]�Y�E����� �x�!���j/�D�U�{Q�;g^��2��j<�q�����d�1�|-�B������iB��
�P���kh~Ϫ�Ԧrk�b��p��·^�[T���$����ӥ5N�P/��~ �>�i�U��P<��Z �y��-��G.E0�����A6i�ҳx�3ܨ��d��sm�+es9���çׂO88κ�a�3��*:�����˧Sr6�T(tUt��۞y��'�F�b�ܶN�5]0铌�h!ۃ���M�Ƃ�*�=��v���i�p<�|%a�k �TP����m( �a�N�*�v^m�Dސʙ -����.��&2QXP[:ȪJ0N9^q��?T�p��\�1�3���Gf�2�\+�83���H�ހJ����&9�����Z�	�`�b{d6�����:Y>��ҿ<�5w�vk��[^����cc,i @~w�)d]�	�|4K�၂�J7�s0p�]��j
��n�<�G=�n,*���{9q������x�Ćׁ�Ȁ=�������I�v�����`�4!19��N���һ�v������t�4
u\d��G�Pse{���9�����+@GG1p�M��؃�v���o��D��ٕK�(�'�q�{Ҕ!/��鮹(���) ܣr��T��a���&!��\<�~I������@D�$b/fz|8��x��7�M0���ݡ����9�y�"Ao��FϤ��u�J�a�1m����V*���\��z�0=r��j��+�O��ͦ=�}�
:�9l�tW���%�ZР�Zb�V:�R헲��>��[�MRO�c�C0L:i��s���W-�u{�J���έO��K�]�n�M�݈�ȸ$[Y*�/�E��Q�p2��s(�n~ԅ�
���]3{h�������Cy<�H�\������fM�2\�370�=��ck�2¯�]ݿ��g0�GBZ�O�r������#Mq)j'��~�����6��)�]��I�G�D�ٳ�y�'M�}?�	� �s/\�2����}�����&1�Z0��ʘ�[X��E|L%�rd�������� �zF8����ʲ1�T3�ۋL�@�j�2q��zu���>D��/�H$���I0l"I��Y��-�d��g(�L1���0uX \�c�f�1�A��i���ز�A!�?*`Z����:�$�`r�	����9�4�B[G#A�e"�Z��e� DYxoq��v>݉X��2g (t:˦��-�A� ��Xf��P$�`�Dr�
���/�=z�����w��G�ѯj���8�cjjY(�~fD&�����t�����/���bB}�՚�u�w��=� -��'N*�K|���&�r�����F��Z�ڼJ�ޓ	(=� ��.�v�f�������4�P���$V���¤�X@'�i�t}�I�����ӫ�C���BM3�B��H#P�0G ���[�_�G9$���2�/�
<w�5,㏾8�'&���u�*G��<.�vcNr��W	����Cc؝�Cy��1Y��Ͳ���*��V���@� 5|�_8P�[�Z�U���1��Q��Kӈ7�[�a�3�bDB�K�ܺ�t/��
���P�$�/�d�,�G��k���?.
�e���1/}ڍK0k�%^�Bn�!��� '�m�%ҍ��m�3{L�k[��k?�{n�{��/�r*�qb��b�c���C���'t6�
����?ꔧl=0�!���(�?�Qsv�b
+���0\��F����o�c(6��P��[��eOm�٬מl@��KZ7��٘���������?��e#\�eL�B�����=��d&�m��p�z�"���7zǔ��Mh��s�{��_.I�R�������{�@mĽv�p��J��j1@;���� q�w�L��#��	�b������mi%�kB�b��0&@6��.AuÛ�Hup�3!��a����ɳ��a�!���%*$P��� ü�&<�w�� �ģ�$�;t4��d꽅���g�&��XW�K�4�g�u�KP\+�3Z�C�͡)���ʲ
�OrD�s�l��6���X��7��0�aS��I<���&�T{�PA��ndwܔs�HN�B�Q��ў.��¶j���\ز�wNUsE�I���&v�KZ[��Ɠ{ h���>�G�w���~%R��ܠU��+��`I�%`~2-�<�Ɔ��qP�zX��&���c|v���~���0�L��@�v��A(s9h��u�˄ �D�P�,)$�[�5��E��i�ETy��M�xZ '�U/a,7�d�[F�;(�����}f$���B{���;9�!�ಘ�����lT��t/�4uH���6(s�zt�8'�/Z�03��x�3�=�a|�a���h
���Xsj�q��V4Q4��NeY�L���.�ٽUۢ�Գ���;R	�)%n.�s$�xG��N4���=y���\��9k�U��LmPO۸�!�����^�,a�kH/s��w~yC�znI�~��հ���ߕ��t��j)��*>�� +�p��(�.�����~d+$�Q�&
�K�`�U���_��"S�씈��L�=mй�a����f�	BDMrUw���ۭTQ&���L7!ܛ�"�O�ع� Ax�F�q�˦���n���L�O�ey���匩G	�p"�}>�F�s�z�x���)@�hWc, ǭ9l|��LH�9-H�t���RW�z<��{hͷ<�~X#�Vud�������kjf7O|ny҅yC�J�We#ӗ�ێ��>��V�0+"�8�"&	��l�R