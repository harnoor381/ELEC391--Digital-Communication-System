��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����,�1	�)��&��(��H����dP7ɨ���:��0����,�6m���Ib� ��JK�yUh^��9���E`���K�
��Q/��V��T�"���-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_d
�t!���N�S��گ/�TNM{�C�5���M��;����L�S�:�{���\p<��)�0W��B�R<Qt��Ԁj,3Ӂ�v��`s�HW��眣�U�Z.͓k���ŏ�^�sGt��P3U����ŷ��T���O�A�LM�-F�0��`86(4R���F����J S�[,�+�ڎ����Q$uꐠ�1,J�l���.j�&!bێ;�8b�أysH��Uˀ� v1��8��VR:
���N�~��$(���l��z���g�1�:��׋` s���LR�$�n�����r�����?�9���*��ln]2n�t�3Kݤ�.�Q���
�j-�ZW��F�GU`4�%���}�4IA��_s
t
��#�3:�)� �cW*�؃ bh�.�dD��hz�Ά�ӢAv�h���� �������h�M�L�����W�XN��%4�^���|ӊ�.T�N��#���"������ّ��N�å����[�yb���E�
��¼��py-��O���SnZ��vb���D�|��Yn�,�!)���No�=���v��Rt��.,ɏ?{��f �nE��:z,W�w�3v�������om�KA��Ga�s4�ƫ�b�t$�gE��U��Bك��JGkĠ�D���FD��_B鹞}�2���v���[#����a`LȖb�������%�p��'�R1��:ߏ_�����8���r��M&�/�����^�V��R��h��T	��@�E��@�����.උ�c�m��nS#���Ӆ��H�a�O\�ų�0�"WK,m� ��J˹J�C�L����/���P��ޭEԜ�s�8�=���VW:`� �N���	yF����iʬۉ�lV�
n�:�tuو/�'n��*��Mtk��daL��G�����E�L|���(����V�{1/>��ࡏԮV
y���C��� �����L1���� V�|��]E�;���@�v�w�E��p�27�}hi�C76}z���k+Ksdb�D���MԢ��wBp��,�U��p�4�V%b��ج�/�iO�未��E�˸�}C����(">@X�ܺY��]�Ѽ[�q�E =!z]�5b9S�*g~��P{CD�D�<�c���Y��B	Q� F/5�/�]!��Vdy�H*�\z��R*껃�4������F��9���7og��挈D����Ȱ��Y�!��1� ҼJ���E�J�3Hri��_~�-����^ް���B�߄EF��;H��Q�k���L7�����̀?GY/��D�:�+g�~�S���"{!���}y��\M�`�cN.����0���d�U���ZtA������,9�*��a1��ܔ�}�ۦ������!�� O���:>iP���ڪ�P�v�i�#XYO]�������ۇ��P�����P�$n+w�?��A�}��� �l�a=���aZ	�)G`f߯Vr��(�]\V���"$���|�5���S��QL��<C�MԹ���!r�{�z�X0�ᑝt�(���RV���P�IKj�������Ru�+|˄�P�kr0�a�څ����J�#z��:~@�)�U!?l�{:��
��X��\!�|V0��
��S6���_��5����ܛJ�A��-w{d�Id'(��(�<jFć��p<̙�Ӡ�8�L ��䈑X��J� ���_�]�P8äEc1N-�sE�buY-���*�ϥ[�M�t�E�aL:���R#h�~qi��!�)�ƅƾ�[ B��;zlP���l�lpv��\����Ȃ��Wc��� V�J�?�0��Ll����W5#������e��0��ׯs ��δ�W
6��� �B��UR�I����89ԍ�l��mi�d�+jha]쏞����J s|�>N�<z��Ț �9|�I�xO���i�_g�Q����`��x��|y8s������LBc,�-ך���]F�"�o�M2�:�W�	�G�(!��"���6?��B$WG1����n�g���z����(\�hG��-�)�D�:�,�� p������I��ct�G`hM��z*Q�*Ci��8�3r�c�Ph�Jbc�hW������c�����oO[��0��������\n\\@���e)_��"'�Flk�_d�8��(ޟ�r����� "���ڑH��7YW30�^�D�?ep 9��d���PjkW��7�{�K~���~�|,Bϰ��.����g�5���x�h�fÄP�q��g+�'[�7"�g���I��!wՇcS��=�I)K��Ț��U�|q:����3{�߭��ʽ��K��Ƶ�}b�C�+�����t�:BҫJ�E���8x�2�0qN���w8-�!z."e`�Nm�����ׅ:.���ܫ�l~X3�����/P��"PM�f��*�A����������I����R`:��"]#|$��穙���?���+e��+=���*�<��|���0�5?ʦ����13���P�Gf�W�p<ږ ,l��1�6"o���3�������>���0�q��s�hyb�1����f���:����ix�'��9���f�Z^5�T��I%��b������9k��i�t�}D>�I"ʯ	]K�?�fZ�F$�dEf��H��58������w�֊*��ӈ�|��rl�{Au5 @S��U"`�[ў�����&1��yu��f�2�<r|�6����� ���e%,�k�`��UTA�������./�>��4�N��@�%�s�i�È�	����*��ı�;�e}��'�NW���枸q!�<���ϧXª��+5yޮbcU��"�8"E,:>(����k�����`��l�\��B [4j�
P&���ƾ
f�_�O��ϱ���fԂe���ks^��ѥp[#��6�<﹂ɹBUg/�Je��m���������A�����b���K���h�o�Xq8���ռͤ��%)-;ħ�L�͙�tb��o�ƻ m�h��� �_���5[�{�E�\��������w/���$�(�B��}�@�B��n5g�a�#s^�	s"d�.����8Sp�r(��]Y����M�7���'�BV�6w�0b'U>��	b1.��y�J�=$�<r���V2�,`�[�׵O�̔���r̍!a����f	2��6 �]�y����E�G��gǁ����'��;S��髠���e!
K��]�l��(!����)�z֔����[<�:����-G���H�'_����� ��è��H��oub��Ω�WD�@�7Cd1D�������t�d�����US�㖟PY�����{�Z�j{]�o/
W�v%i\>����N����~� \=�L����7,��ͺp�b<����h'��:(+1B��̠ɔ�|P0x����g
T��ɟ	���U��zݗ�՚2=��7C�4 ;=Wye3�4����q�j4��-ר��u8��j�Ӄ��c3�gX3� �0�U���E�y�.�}�鿓�"؇��g�U��ov�u�L��UO�Fu�B(��`��,�A
=J���I����ʎY��/Y�]i��X�p���F�^h8_���_��˚�P�ğMl��b3
����u����r�<�zП2�O�saW����i��*��%�~W������{�.Ƿ�l6h*�������E!x��?Q�!̝�i��8&��p=�D
��Y�����=�Y��$����P�[���I�7�xm�u���m�ەݠޥig�N�B:��;p'�Q*��9<>���^k��]��^F�b�0�)o>xP6aBYt��\��&�`�%�e6��P�H���h�G<�/	��/�� ����>�q/�q,���r$q�P�,T>������� x�=�귔��9xR��dwu,_b���K@��ꚦ?JA��uN��w�n���ߞ�ۼ�������/W��M0�iG!��;�AJ��S��0$/�Z����ˇ��G���e��κ(�� ��Μ��9�����?4H��6(qn~��^�8� #�����l���2����^<]��ح|��&�R�E�c����C�!��U�29:�z�-�h�bԿfee�t�W-�Xu����%�Qڶ$��Yx7��n��\9��
�狏=oQY�k�&�C0��Z�b��9⿭��(CfA_�����t�ޥu�>������ޖ���F@#�s�xr���J�)��r55ǣ�G)�\���n�⠍���\�m�Ӌ��+A�nKg�m�@�m}��[H��YE�ܯH���"+�&��U>���{�'H��@t�,��$�;Y:��އd�aV��5��X����C.��ʊ�A�&�2'�D?n6A�/˜�Lqȟ��{��#&�\a�_L��)���³;�ҳ����Ӄ �"��-���|�B��cg�<"w��X�����E�ΐ�C���*��rѽ�01ޕ�%��H��r߫��nؒdR����^0���)M����$�q�bq|^!b�`�Qeap�^8�	nC�Aс�2���}*4�$��C(��W���9:���(F�u�F�g�F�k���h-9�*`j�n�4����(��
4�p�6�NG��L��/X�|�Y��L���&9ȯ��(�ÆC���]�E
�$�=���۲��o+2���R3��Q=)]Q�� �9�O'��neѐN�*��R�"Š���6� t��,G�i�&"���T�z��YHO@�u���DI�{od������~�C�&�<�f�?�OJi�t�d��zI�!���j����swr�677����k'@�;�$���ܓɇѰ�i�ov��*���c�����K��&��#�k"������qJvN��h�U�.H�N��)�Ja3�lp���@�8Q	���G�*!���guz�8��-R��#� .�����Z#�bS���a�߼��3��X���m6��$�a�;kp)�s]����p�Y��L��?�m� ��+Z%�Wܿā��T~�Ni����ã��	!�/�^s�z����W�����)Sۙ����"�@rf��|(^�u�,�f���AX�6;�iN���!q�s#�@�5k~�����Yظ+��z��g�n0�m����̦q�J\�o�39�ѫ�ȾU��%��j���ݍɻN�?��3�H��q\�ω������\�.�����9b�
�&��O��l�!e�4X��WY�MlӺ��s>���d;n� ��f:� �hevհӿ�Kp1�����3��;@Qj��I.p��%��kr�#��S�Cy��l��ܾ�bm������	��Nl�=���-���IZZ��I��o�5��G���s� =�Bi�C�_&�<���@Ȯ�F��_�]�З��a����bX4��6E?ߏ-�v
R�~�}X��^v�g���>?�o%�sq���%O�+�"KTc��'����f�~
�=W�Ǖۯ��&���˃�aj@`F�u�lJx�O�ԬG"Q]:��D�o����8�mH�$eu�:���R����0��c��E�����/��w>�D>�$�;)�Y}�u@��MO�̔��%rR8[�����4C�v9O����T�p��o"�rt�աt�l�������ߚ	ⷱ
P��D��R�<�+!8�Y�CR��-2_��.�<,�}:��em�+Ţ�E��Lۤ�Ͼ�� �K�ʚMv7[��z��ϸR�N��)4���W.�����<�(	,	O��,�Cֶ��OV�O(�aC~,�Ñ���A�Ո$"Z�Nܬ�x�|�Y�2�K��JQR��� �����;|֐a���+Lv����>U�q1;6�͡��Α,�����}�v��jQ�i�oQ�U�V�(S�gJB(�*��c!P��lu=��W�Y
@"U��L�0/x�>��~s�)��-M����/!�|[r�VgJ����P��9�xV=��L�AR�吊$a<<H�S����fc3���:��Dp���SLe\���p�78����˖E�'�Ć�$�t�pqZ���RsHԤ�j���n���'tM3�$�Ġw [h�Q����+��78>�^̠3�~E��Z	N*����x{���j.+O��zr�|�~��ͦ��@tV�w��>"o�G�����oZ0�^l�5�"�#)�O�8Uo�鍅��g��ќ�w��_�N�jzU�����;�~�����IW�M��K��ir@ ;x��$kK6Yߨ��OtߣcC�#��OM�s��ٛ`g��-ѷ���C��?<M!O�h��ƥ���� ~-x1H��C�?�f�/��8�}OS��6�2�L�����ݮ�>H%H W�%㑄�P��G�hLS|��j�#������ksy;o�o��$��V�R@f��TZA������NI��z�zXR`��- �Um V36�%	M��K˿�W�!�Ы��./bm��ٟ7d񁝨�h�vC��S�h�Pʊ���F!1Ӏqn�q(�잵�A{�q���1[�2͗�-U���P�z����iY$��y��yn҄�? ��B���f2�_�"�<��]�o3/6�ʀ�L2��Ӭ�ф��'�
�W�|�0�<�%��M7�m6��qG5��9Ӧk��T��x�\C���]�8K��0�!�����Ь��).P�yY����cA��si��$A���o!L�0U�e~x�hq�&�j)8 d5�-ޖ^C2�n�zfL�Zo��r�o�q\���3�,�.W[�k �5��i����Mf�zA傞� ����E��~�A��q��)f��U�)��3�xn�ډ	�y�㵜�~Fh���xo���\êBz���@�*�t�=��鋡$=��W���A9��~DEů�Y�P�l��c�[9i���I��J�=#�f7C��,��i�+z�3��)q��<`_�^{�=�PV9��K�T�:���"���B�m��&'�)w���
�9�P=!L�*��2^���􎠳�nz��mO��#�1��~m���kk�+��d^� �D�s4C\�aR�]-��@��l��i��۩y;���_ui�r������0Ne�C�Н�;�z󈖒��>kĚ�v��Zb�!![�D���,�Q���ʬ�p�(���1?|��Yܘ_ʨcny?�m7o�YNX��{D��.��A����P�\8Oy�T·�S�A��-�"~v�=���XT ���1�V� �E8�'�{���lcr�Q|*�搜.�(4%Ҽ'9��
�q����k{4�|cs�s���e����4�cY��x��k3t��Q�.��>�k���8;��zEi��n^=�� 8:����I�X,P�$�����=��l�q��N|��0#'ڃ߷ 6$0�$�5O�rQ#��8[u�*�<��s�з�{�,�=�-�s�`Wa�>2NXxg ��M���{�K�u����-������P���Q�8��U=�a��/��##��5]m�����ڧ�L�"��7iR�>óA�\k��BYHhPJ$8��v�����w���^��4;����u�Ab�ԇbu
ҙ��<��߰�!�*�sԏa�0�k?O��Ƽ%9Q}���M��G��
;UY��w�Mպ�9L�F��T3�����m���S??΄�g�A���(�����@��4O�zx�r�E�*����?Wjx�KEE�j��O�˟�J\��*BV).�BU�3 :0��!]��'�#�����y���e�H@��q�ϫO� �xw�^�|��ɫ�������`Ɲ}���H��#�
�=E��o?���gz��k�i��a�ɿ���u�vX���v��>F�h�j�9"��`Lr�d�z9X�L�����d�|��י�ZI`��7���:27���P2��r���B�GeX�v��E�l ��������\��QL����v��s7"�L��]hr�84#��vA�G�ԍonEq��yՇ�w)��(pK��5;?Ͻ�1t��T���Z�v����p>؟{)W��a2���ty樺���H%�ڀ`���H���`(��hL)H=��(������U3
sz$�݌=��';ރL��hU���m	�˓��BL�.u�ɥZ i�H6ŨPR�v��1�'�>��P�lKK�+ \�p�5`��E����dq][%AN�y/(�;c����|٭�Ht@WT���_��y'ü��-\J*�2��y��WǶp6/0�&%8�T���䖓��,�wT0�=A�X�s M���P�:��n�w��Y.r ��"�������ĺ-!����=��ӻ���[�W����\�5�������g�g�񀞁]�o-��%���U�6�TQ�&B�t��I/̢a305�m.Q��Y��#����dCn$��Q>b$E܍����9o&Ú��'���?d�Q�j�&`�^�F�m>�#.}*FJ4�|=���Y�!���
�Q�(�)�	a9uo#�f.��l�6�`���L`d��(᥄�n���U��ؐSI�ý�%��СBY�ΐ�F
(T��I�3f����`H�n� ���:B=�����|� �6O�����4�UCj�r\h��i�>e:8�a�-}GIf�kq��L�J�U�t3/ߏ����@�)���>r*��Ҡ��H2y]��Tb>L�FK�h�}Eڜm�N���}����e��|�f��~�<��Ŏ�e<���8�4��-P��5��+�	8��";�^����5Ĳ$��'Z7a*��L�]��8�g}1����?�E�4�F�kS��nm+x��DF%j�X"U�_l	.�����R����3���� �޸�� �y��aA�Zp���0�m�EC͂+������;ղ���V���;BA5T�S��m<�����77W;�T!J%����{���
�<���od���S��4Zm�].�9�6Ԡ[$bƦ����#"�ˮZ��p��&�3̥�(LT�H��`qI:���W��6����׬���X�|kY\�E2ps�Z1P�vÉB�6���Ξ@v�$`�z��i�V�"� ������A4Fųҙ�h��9zWY�@4�;���F6�Ī�W�o��gɲ�0����x�ݑ���[��f��'��eV���Lqn�3;��M��Z��f�7��)����RCL�e�+/��[d�l�\	��2�Y�����A�\��2{wlA�N��H�҂�aۓ��Z2�mNC��[�b$�/���+`̓V9'��@�J:�s�0����U�8��5���n�j��OƳo�

�m�\⸀1�U>�#	��Eھ�#q�����!�vT�l��vt��C�����Qެ`�D���3:H5/_kY�dv�z�8����$�u|�j�*��j��y��}��8!T�U��X�0��-�������1:(���C{���EG͜�M�^��qk""x����{ p����ɽ��� X�Ȫ.��'1l�Z���Y�-"X-���n+��q0�����%ߍA��P:8���4^=��')�D����Ă���%�O������8ý�x��n�HnsJ[�E(�9��V҇��o���%pS*a�)��jC�H�׎����Y�S�呥6C��*��"�[��0��|OS�:�4��2>Ϙ?���&%6�4�d�1n~O�D�� g�ܳ+>���G� y��u�v���Y�s���0��[Ȼ�&!��/�cސ��/z�J�wĠT0�Z,�_�ME��JE��=�ă�#���K� �L�H����Б�G=��}A�P/��MK |�:�7���/>�������?���RŽ�T�j�h�w�����"/���pdaO����FD}!��DH�=Q��s4qs��6]��3D~A��(�
�-����������3�YG��ػ>��0��P��8H܌�\����9h��C��a~Y���b�m��ZaZU���XZ�6&���ʀo�@p�0~ːC�.��}c�\��(B��P��mκ��v��������H\��T<k�t@.%**���n5$���­
��(o#>�c�s����i8/�Fq�4B�� g�[��Q�E�.f����.�+������.�4L�f�5��`U������E�Y��_���1�cIE:�q}w-]n(�n ����$5��sv�d⧣���sc���Ҙٸ��fhRZ�T|*����昧�󭲎 �M	!ڪh�XlE�<s|��r0j1p�Z��b��	����Su:����>:�i�i�$ߩ���T'2$d��z��#7�JK���
yү�x��tɰ���8�s����yZ��I4𢣉&����5N�}��#�>YW��JrDb����mhą[�~�Tr�$���`r�5bB�φ\�k�(�Uw�0��V�ҙ���� [q�.
~O�uN{���z?�̓��N��J)���M>�XXIsYF�w.���l��=��(E��I�2<�*���7q��(G��9b��'54ȿB���
մ���uU	nX�}Y/l�������:�5_�� ���J�׀-�ôz�`��~>lm�RԈ�)�6S���e��P���\q f��y)���A��Pg�~�q�1F�gٻ������\|��^?H���ه(<����V�:Vw�����9|�h��=Ѥ���h�.�\�Г�0�)����D+5�K_���>��@t�O��W;�P{�v\\�q������H9�����
�7����(;��-j�<��G�8�;�|E��$爤���F��M����ϊU��wە�7$��ѭ)�N
f�ۿj��5���'*$nPp֒J��*�^�X>bޤ3�Z���$��Mk�kH��f��T����g����.�pR�9u3��h�5��7�� �B��.�Ot68��G�=ϵ����X+�J�0��dY�o<;֍ ��1��L<��Ъ:�>H��)�it	�	M�������4�B��)E���D3�)lV���
mp�W��to��k�Fн�{��!�}G�p��bΝ3�V��jl]K&^fxS���%�V�P�V{���gm���v�n�uZ��?b.j�6ޅ�����&������'�K� �[^r�Z�;�����ץ5]� k��z� Jc�\M�h�o�Y�e��3�hr�*Y����O�ѥ1C3���������骢�4�4����� p�L��.��ݸʝ����U3���I�G�p�[
�G�Ug�mY],�JZ)��E�x �^SGz�@��?ֽ=��;6O1��D��* ��'KLu�aklK�j�3��IF{m�o�]hژ8O�B6��{/�u-���.o�̢ �x� v��Sx1�<�Yn��%u�X���}��QG���w�-�	I��M͵�+�����ϭ�^�^�:��g�'`����b��Z��p���s���k2j^��L��i���3����[�#c6G{Д9h1'Z�-Hx�A�Z�:g�3�����C�\v��5Ǖu,��`B����6��P���G؝�iN��FQPI���\�m�^�2��;n�U��U΀V�*n�V�� �Ŵܜ��g]��=>���Z9�PNH%S�MRW~�?�!�D�jS�Q�A3HfV2YO4�����<0t��c��7(2����B�C����c���*��b��֘�l|6�
��\�ANՅ�ʛ��M�L@:y�r�j�5W.}tQ��'�f.,�e�&'ws��K?W��[��\Q`:/Oc�eF̐"�E� �y��NcH�,*&JZ��������k�f�Ka���C�q��#��>�g֙үBQ��zٴ�a�v��@�0�)����N��A�C���HP# �U��{�H�����XmN��h-��w@�Kn��h:{�_�(kS{���Gx�}��!h�ݻ|.T��d�8�v6�!ƅiswFH����b����9[���Zu��㋕����Js����RC~��B��J�B�����S�mҧ�b�e�"�����e��VAh����$�T�[��Ѕ�j�tW�x�8H���]2nl��y��W�tQ��zJɔYI	�vd.j�@��~4~�����n�j)�	��O��y@7AMT�}��Z����E�3��w>�p��8�Pu/��Q����r�|���{:��ud��w���t�����u�^}��*b-y�x_,�g��^_ҟ��ƷB�1��s
>k����]���q�����'国U�A�c��۸w�*m�&h�Md5F����:9��\��T���0?�7� �d��8�GiU?hцl��
��PՐTP/}�ɞ�����o@?����Q�Xp��mA�v���}k2ݽ���J������yY�uѬ(�U(��En�%(ʧ�S
X�����|���s��	=�3 i�ŀ�)X�M�?&.�����N䦖�K�T���p����ė�T������@b�?{#���/F��v�i��0����S2/(�jm��~�ӐR%;�p�\O�9j��H#Ɋ�&p��~�qdC0A�a _���8�g��.���Z�ؔ+ׅN^�نPk`�I�M�&�������G�}�#���"E+���g�k�nYiEy&Je|?s�HU���'����*8Bg(b��������I��Hz�\�{B�8�F
�չF�%�2��0���`�B���nnj%�^�l-ӈ��\�U���h�����؝����;C
���9��G����/�B��9r�Z"ݭ6*�$�@]sf,7�#�Q똦�
�����3r��Ȭ�?�`�?�eDmݧNV�q�&�%1��8Tj��5�y,T~8;[^gLB[�.8��Ӹ���4���<~�ʜ���_e)�_B*+��S���h���AI#�]�u���4j�B��@˥'(��ؔs�����v�$����X�Ijí�n�����3��mg�Ъ�}ʂ�i����//4A�������t�D���Ǝ�laK1��f��
��7�	ƚƢ�\m^�}���C�i���Ɯ)DE=�������\���Td��/b��:�I��fv�tny����3.����΋YJ�5�ںE��[@q��3x�̀����f�3�Jְ&������l��;���@���x ��,��	ډd�BS~�@ ��������ơ���D#V�Q/����`.���+�?�v��Eki5c?z'���?��$�isT��U�2������������õECk�朩Lo؇��p�G��2�	�q��p�y��i�U�VF�\�;ѱ�C.�"�X*7!m*WT�)�����ɛ�J� � �/�����L���,����#(���ArF�|P����A����ıf.�h	!��R���܉�up�yD��QOZx� �ܵ2�y6�(H�����!�F�n�c��/t��e^���;8"�(OO�n��Kݬ��U|
$ ��[��0 �����"6A�,�pz\��|k�AO n{�"�g�t��
���K��C�������A>/@��bsi��6����UM��{36��oI1�y�Y�V���\�+6سBvƯBQR$m�H��-�6Ƌj�Ԥ)��3l��T�ئ:XG��G'�At�Ɏ��X�\��׃K+�H��z��$/+�h����=߷�G(=|����^z�2�������x�E4��0�GY�62���gl Z�I2�8���a�u�Qv�_�@~ �rV.�j���l^�����Rn�E|w��$b��k#o����5r���;Yز��l��n�t����~�p�R'b����V����8��7��� 9>�o	�&��Qd�%{[����R�����N@���>���ˁ��bH�F�B[j�brK6TȊr��-3�0����Kn�.�#�φ�������1�Z�� z�:��s�$BA��Km�0���	s==�f�q�58�`� $�����&�
�Ρ��*��Nm�8Pc���v�]Ձ|�Jn�y]a)�[�(�7	Ix4��Ouf�w��bn�"�EK']�O R�kq3歨��z7�����רg�Brp��;`��'*e���R��`�)�>���E_N�*�8�y�T4�A>��!� �+&�K�GR��a��$���
�4�?��zğo�e��|O[3n��Ѝ��;y�����4�P��2�

�r��3͠�5�����l+I�����HA����ָ	!<*"����$x����� �v;�q����6��J)q�
5g����s�̥p�c6���2�$���k���
�iz�A�	;AP�+
!�.#`�%���/5�]�ex��yqqٮ꼪��N?�V�46�5b���r��F�	V�K���I��鳷�tx̚�#�����J+����<X�-�)���'�k��.|7���g�#�Rp^�jӼ��mKAC��xk�8b�7�H� ;�c+t����"U]�֤L�̇�}���a~�NU!���8�F6h�N������Wբ�(-a�&�FN��$V�l&8)� ���\�ਈ�N���t�#h��0�2�\_��fz��AFP�h��c��Xkn)����4�Ԗ�Vc�ӻ����`�|'�P�y���A
n��-ʖ/�L�����oE�w�vl=�D)u5Ȩ|^-F�35-�H�A��E� "�>�Ab��ɒ�yL[�X4y�IC����'H��H>�ʮF�X�0�D/�M�"(��'�~z�x�Gs��+⇎����',�t�6F��f�[���h��ۨ��NȦ�e�T�0g�� S�'�U�?_�~��8�D�jt,f �%{e�sP��2�
�gv[�&��r���6�l9֟�Z���Sk����<�K;��U{�h��	h��2).�C+�aR��J�^DU�ul,�R��XTe�1:�u�!�JA����UA�x�U � �^�Q�{z݀lwd!������蝟�@��a�;}��	����|���j�l�5��6��9��h��Y�Y�^��H�}S�J���G�G]J�KY e9����y8�g=�+| �����ձ�0*�qid���E�Ԓ����:d�7Rg9�W���P!a~/�(:��t���
N�Р7<,�b���%c*�+[- �Y��݌�c_����2I zVY߹_B@�����M���%R�:�����C,�\�J��vOYzT�j���Z`��d�̋�2^%;Jζ��Fzp�d~�K�Qg�\�R�=�-�Q"�cWB�;�"m� \�S�@v�Y�%�n ͈c�C�\g�0q�V�l�FV���E�l�Y�N����P'}�L���]N/��R]_�K
͑�nћz���qsz�qM�y"h������Jd>q��y"��B"���&���Ē1}�������x�kPA�O|��V���`�U����
��<z �����S����^$��u"�,֭-�x����[���|'�����ě��f���N��h��
?#�P�#샕q������QP�|��<=h3g(Ĕ�����}�.t�+ັz7+G���u��8
�,I�������d���g.��<��w'?�D��"��fZ`��N����A��ƜP5��ns�̺�P�R�xJ�䣾���b��uS+�
���,D�S��}���Ջ�R�~������3mk�V�sCј��*��m�]����A��M ����M[���CA��������mk�CKŵ	_bc�+I�aW�D��V~o,�z�ɤr;��)� S��U�O`I.�r��RA��ѭ�x�b!(�y���.Ȧ��"?�WZB�w���7�"EL�~;J��J�ڵ���h�e���AJ~���s�$�/e�%� �n��T�
��
ب�1/���$-<M)ϭ����b+/y�Yϵ��Aj!�i����2��vr�a�*1�