-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
gG4qAjS1FmF90ZdqDlq+t8nTlvXZQpj6+XyPMVxWvv0m1yNAWi2QNg9r3cV02QpamVcVpYcSoanD
HOYt4ZDfQHwNYFyn7kikvhhw7NeEFRZqliJK6N9oSzj4+3vQLz2vIYYuRm4IoJaA3aq9Sd3bn7fj
tLjcECQMJddalPgALf1pwre293Wl1NZZkGf+UZs/LDymZLte49MCkMLgtHBPmqumozRyJh9wlTJt
6YK7aXhKMYMs4u3qqid8gwNIOIVbilZNW2yLNV8JrPdBHmoFc68MLzphmKPWmdNbk76GyU5uMnWL
JmZetUnKPVn8Krkujkh14ixwrpIR6t0auxtzgw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 12688)
`protect data_block
2ApN7Ro6lMqIck2Ful6Zn+gR0JmCa3wDEZ6DUn+HUqyqTtndC+gEvahtZmie/kmsk0EWHOjezFsA
4Ej6ArkNNDxfI6+or1/brwrIs9YOkbsslion3hAap5TY3qAOS61PbOdLtfDdisJe6jiUZKh1Ohlg
kGpswRk+SxYYrXbQu1COit4S25LUvA692hoG7eo7llmIK9SGH4L+7HhNeyZqdOycZiOqQDHpnKiB
FmZ1diPvqpudMeAFGSDbHsJ+B50Mp/t3JsFHCMkqU22cJbALFW/KH3T0g3q1UzW2SIhHH1WPu/x4
ig2IY2pIJDSxLXAWrCJpOLhMIH3NvCkOFAzaUyw6mtCZb9m3SsStJVPJ5dlqAcgV4qNQ9gCPicPs
PTAVrW4pELYCB4D/u8RRRvKPFBdI+3g5Cu29aINUkGERlGx6FS/nLDyM6sLosYUGTecBgJBvPRlP
bgAUYFzPcGs7pKM1JiOBR6FljfLSo5J7+z8T2g5eDAMIDFBjWOkMIvsChCEqI55XSQN1LmlhjjhN
hrHeI7Kw4NEDi++aQliSnvP69HlkDzK52oVJhJi2MsKMwvDTVL6BIGbX4Ma9axdTmautU2PI+OIN
JMVpzs6oqJX8gDYPXouB0Iljs5JK54jCuJ0FAHF6k2/Gz1uvY8MJLOrVYa/bEYaLEAVKtEWEXrL1
gCxyPgnWjes5ZJCZatoeIdJt7dgeUqkCyJLkX3j69yt0OH2zjnqmZ3B5k6UhTpl4HBbuRZrK+71T
davCxEytP0y55J9lFwnxMqrL8C7NIg2nTZQ4NMwYnh39Z22dcLIPrEVRK33WlsJ/zmyLFpeW2SVX
LFjZ7vphTeQzE8btwEdAeHG5L/kIEOl7/T0IzilUbg4OvWxXiP0i3ovS+gMypGPis/6n/n1MzJ+n
a9+ZQ6yyfvI9DtXuHbzQrqiX6+sn5C6pNJ0ulqFFBBQMLp4bZf80eRe3rdFOdWrMqkAJjvex2pcr
clpU48FL6qIqUnqy2HVDiiSbR7YwqRQ2/MN4m8BGX1PdY5h2zJzKToWv5pmErJzzvCzM1VODedMb
aFyVm6rRUPMBpF7QJNZaRZiUHFZi17FqGRRXDdjvEA2FSDn3ep4rQT43sson3RU4QJMYao/tID0S
B+NlNiGJqAGdZ22n3S4B3paA0+GpU61iyekeezpn/Qr+nNcuNUSy+WKgWvpYUkcZmmAhCTIl9Kvx
hfws4HjPpNMjsWjhCxGuCCeMmshgvxNxjXeNmV0X4E2x8ALD/ftR7TMeOs0Z+tMiOQamDI2dSJO2
BHngC1qyp6Hzvf2PlJgc3+Dnb52+BA+lO+wUfY9NLVzEodL52vP7nBc9X0DdYpr/uWL2qWws6x8/
BZkv7bn+roNODnsOV9kfpMBFgdAYTa2Pwd54lJvp1vGLiSnWfYhkEvjC118yOUbEkSagJoaaxOgU
GGJENOZq1zAYCVOoaZWuxvB4aP+EsW1p9DwJphGh4wo8gUaIxCCWKLq/B9IA+hWbi1VCY5WjY6FB
UuiWAXPqMrMUIXp8J51WY8NS/SZz/2Sg2ZzVZGw0HCKu8P8eAdFoqeRIczYGkX47NbYPCi7kI7Uz
0nBGQkNrS8XEKq/Ivd/3vs6f474u8ZzRVOG9F/7kEmF3Lfk2ly8MOxBFQgohyuW/6wtltXgklwsw
AML7/cHrpuF8+OMnx9J7HNOaLlPF/VQyoGlpUGJdqyXFNKTdN4kmau1KOywSOVc6izmDSajfH0+8
P3Novk7w2YrrVEOPV7TZvx/DIPcjRiQialfMuuX65pPjoUDpABoU50bUuzc46u5lYmVtBn1E4YiV
hl5JseKLdoGr5+RHX7eFoh3d8+nC4At9I7Bfl8XP8spK2v0nSTHuT7bQhdC4bdYPzClJV78dtunk
qO2u1b1ke6RvM9Kz4Z4qNsFes6gxje+Ktp+L8hhRj9BWNN8SBp8BjYnK2+1Y1WYIniIsBpyfBZ/P
O37GSy82mzC/mhPj37+gL+BH0qPTVH5Thv+I0ZedB5AUNLnJslHQbIFuOMaSXt5kDc8ENZVobNrs
ew0+5bM3yKDqStrwWB5xWdTNYBZOrAeYNvlgP2+ZJgSMbhzNA0h7empM3D4kptX7XpXxWJED2ckU
xKba1cuBd+Y3LWKSeYcUFdkWATx6qao+7991X2yY66GkUQfKmcHm3OwZV34RqZ6v6rdfX5j8zZsS
GLX8/yGHWJiG42qcs+iJTeDbsQaO1ummugNXNojn1NFTQ7PlLVg5vU04I8pe4j8733IIla8UF8SN
t+sI08W4xRvSOaueAzVvRPUBR8ypHXQkNpBLsu+4T/mPhfx9Zqpf+xqBIiLKQKKRR1miWremIw9C
VOWb5Jwj1HEXjbVKLCjiP6AwqKUPD/FxVSUMF9K2wCT94Bu3Ay9pvI9BnQp5fT6xn65kLqoNssV2
70yjRDGixHpnQH2c6ILwCNcqMHVtedpQyThS984p97UGUuuGkh89fyyQDuMmqwWdKCehf3Q9rGtP
7ze0j0BxqYtuZFd8rFSFy3E9TMFJwd6ftEOHQUviYihnXOn3o3hQypFcJBt9rWmZlBC0ykbn3y0h
nsbLjjiiqFcm30aGudfd759nSwOcWq3jAOu7yaqewhrOYVtvUkpZqnr92MPaPoqPhDy/FNvotkTX
tCF+2KG8ZAAhLnoS+xi5rO+LFF/2yiYx1Se68DkVnN9K99wCZuwBfhw0aHPcGOHal+HN7nGV62Sb
FGkQTuG25kjYTrQoYCCrjHJOURb/cwC8ldy1zdWFS0+7wCfKx1B3HUWaef1QdxmPq1HSdZh7TTMQ
5Ri6vTJvpcWQ4Qc+2xczApvq8wI24irxCXdwSZYLkfwFmFZPGRD0u3ApVBpnTPWORJ2Tn9RV+R3f
jYOJtOjVMI9TT+AWU8CP/0qEzhelYznViid0djDv4HKSIN99iVcs1vrRjaSywNrVP/21j5XnFcmw
Mb+hAXX+1zT1sqcmpdGHinGnc1Q6z0HQYe5fMSBTUYa9C7W/wpH0yeO2/u6wMrYdOlGrOekVPCXg
1p6NKm3DQcgebm38FrkYCDBKPkoEZP2ezXnjt1hMcC9+E0qI7cFL96sFTzxLsaLwzOjfcPiPQn44
KjnUt74a2zy/VGdYPOKMf2OnXiMoST64WSs+uoqRUmii4gVdxQnpQktt2fRw41EpX2WEqLNnLO9k
KSvGTpq20g0N/V8cU6nRmgtyB+ZEIt/Rw/Jth4QR9nRJnznvmWIB/J59iAK1knQMQar8nGMUvbZ2
/tF8+2+q4SaRWCV4WKlnvfFMT7dXKY9E4nQtcYFAciYHX1Ei3Fsjx73rxvf1Ld2y6NNXhqDKoC6k
4Yzy7XkqAVZOAEfTpnXsE7eQttCRPSeyO+eIjJuqbZ1212aNQMlFhGGbjFJptEP2BbOZwXdKUdHB
BzAS7gTm6BIbVIVk3Y0liWGf2tvkkM08kLH495fYt/wBanUDIhWSc3EvdWfb5mpSmOw5XDPQvOoV
dI63y+i8rNc4x5JKvjGnNHyl2BPmbVeQi70yoqSKRMBKjGme4syrVG590bmEho2FtdvbMxorNKCE
FUbq4j3X13b18NVtWysJNsYUMZmcnzuwhIe+8PFi+4BzqrAQeaymZkkF/ICYmGVrdqbXmqbE6cD/
oMP4AGcTQ2PmGK6E5LyBVYbStvHRJP4DWfuT1s2ylJlZM7QkxNY8sZfwCcOBj4W9GpxFQrgoRdNH
gdsZIdsr6Aa091IJAotwSsssY3Od0BWqgedBX9AKieFvmZqoN760+4XE1kcTR7CBqGXSG1LK6qQX
Dfz2g8bN6qH4Ci3Kk9Q629CZK1Iu2TNz5e1Foheg6zRBY5n2aO3kQHAfo2CSQPIyM+o11/6TlBbR
UIx5BX9/by46vcKGEx6anXf7GqC9W3udOVqNr3GmYrgFSrJyarz7AZK+NAFE6DWOZ0ZEyBsUROw+
dO4iw782ETbABiGtL1jO7gy+lYStITQbnnpTsw0pvOevj+g92eTtoV29RmwyWzJ3TCYOTwq3Gzh6
3ntW8TKl1j3nH4Xam8AtfRNZCu/gzAd1gzc7an0dIXmbLf9FD80cKrH+kJVlvTP7AqBEeqvDc0xQ
TqgTx2u0PLiUs59GCOYP5CIh+leFL95ZNFqLJrNt4rJUOEDIyE2z/uEz8dEhqQYjrKWXncvNGsOU
LH0JDLpTaL1SIQqCtuEvlTDN+0SKWLHGwgN5u6FTSbBEKv0sitoLOtYFutSU5pqd7t7OIKIZzPJT
wdERgSPuUhHqvDEaXT+7/EcaZWXNZa9W3+ZnAr01LqBEH/Uhu/vUe4m940TgMQwe6mPq1fuupsOP
Cedte+qnAgrTuPLsstqKXPO1DoOgRiYlZedYJZ4ZHcfQjEt2ICEgZo9Lku9EzOq73Vw9ThKKsMmw
W19BJ660H19oGdp7z1ZRwso/Pe2zSt/245x2sdZrXoopMClXqFdFn7AaRVwnTDbGK87VaUYw/Fcc
+sia2AFUD1OicYcbBa1K9DUjRXp+DKng8V+Yva19Xosiwey6G/ywq2OG/fV1a+XW2ELYRY+3u4V8
yiu3PArJSJeeTSLUJRWaignklVsuEs6tUICRH3W45Osi3ir6+9mRa7yZZ5FZquh/K0hGNRl/0xWU
kCCSdzBNDcQWpMOkxRpb6nTgYwlkZP1/UQI9YjMSiqoScepBEmKeHX3+12+n+dqx5xwRhadDAaFN
xShf5Fz5cwx9nHdi+3V2Mt4nQZL1W6hJqhgZurTo+oJPqXhswe7rahPXGlllwe/dBNfOvbA7KAtC
GKbD7Vui6ZJ6ymmoXQLzslrU2mpzz0s7sp4OPOM7vse2FV8ivQ1U9Ovh/cJSQWPhXLhqZ0EiDIvu
CtkuhKLCdWZNIwRTNW1VQcDtCK9AA3Bez+CUE7VztOTkwO30+Sut0ZmUSPbykxsPaj31vXi/uUmo
lruoWOhm8vjQK6aggEjXQXn+Gtx7fmUH/Ewpgr6IYjXBN8bFfvipaWkJugKYKOxBdVUJ/MFhh3/x
SvexJ/zjsMUPVvK0OxdtrHrx1/QolQNcttOEGqIVhKf26jjfzTuuoELM383npYZcIgQ9NWEqpRL6
BAozRQ3inzlNN613rAAxllJqScaiLW04KnNwlctRCfllD8Jgjli0RhGn/x1F4fRmab58okKpBTxX
YUoNT5p6oP1yu6Wy9CH8FcDALYb2SRcJTbUQDuh9a1ijxRNE3PnrSpuAMg/UgXMter9srwgozCss
1jpBasyj3OwGmeNjqMSEdxeNAUi2GdqGc92guwhQi6PJ27Z+II05yoKgtg3QFK/hrIvIGmrndBcj
OVh9NlReFn09FK8VJlL5K7+vlxBts8rzKQ8ZdsZxb0JPLZ9vNL0pDHxNj5yhNY99ubj2GzgwwwQt
ZRD03RwanftZmgJE9xyeda0lJDI4Vn//REG1mhSlgzRGBEaozN3CEwQD/eheMAljqBUbW0ifS4N0
GX7Y5tVDFAhw3kqaY5WfeP1BqBkJkcWV0SqSs/a3pTbBhxU8sILRcs3e4+hGHk2Ci/NVvw3gH2kS
9nji6AAsGBF+zpNOw6MY22rk3+aHXZFu3R088b9BuI/AwhWvmQ1oBzBsN18Hjyk0Jk7wXz52YJOy
o5del4+lEUtGG6Zdgocui+4ph865/VxTK/7NwASy+ZGa10c6Gxf1qTeIippEzrEUfJ8rgiOS656U
1S6+q/nLiNLYTJwSLd2YgBfmuhSCanvy1x45qXvy93F3Tf2Reabec8Tbppep7JCQUzWHBkfLwxdt
Ku2FjtPs5ibgY9Kay+qfiUXnp5T7/2eGO/ua8HGgNtUf4PVianhlzWKn6esiQsygOflXdK0P6CKR
b74LPzALy/f1uMjdE22AoXITMIsjmDjgWp+QVU8zK5t0nHTanvOh0lgdpImQmS+/laQ7n9pD1x/W
YCKfrKB3canL3eMU06GB+EV84e+KyWT0ngwn+OuhlqnngqaNgAZeh258+0GPFbDwib1fxLXprV3U
tt4haAHvjEWQJQWT77Fwj/OI5XoCBH09zHuastvR7iFnNuT9YBcbMfyUE4Sfv1/yaEXa9CtHlX0v
ZRxWrm0WtCcMiXCORTrAfem2xsDTqZE/9twYC+Qvq5IIWmghyKnq6A+2uLGjZfMy367/UjZ8aViS
+/4f1G0GUko2WK3LjNP6H5UsUFSsVfLikEbcn8e1bFqADVHT9oJz8o+tUJ1Bs/mjzBqXB8wBTZVf
8Fj9g1W9YpCAV5nh1YpoJGexL+uNSj27V74LLuKme8QNf258wtqKneX71Z5mNMBOkxjqlBGMPFo8
O608onhx9coqjbwWGOiarRRUX5dyO0IxSMHGKuh7bHVhyWZXpy+lfO1CO7UrvzR0ALwzOU2p4349
Ah+PDbygTgF/wFkib7jDgRLtRRyBlTzlO6elWZOXYtXCZcwyi9UeLT15sK+hcooBjjba4Z/n/X8v
BShj1ur6Awy1gcD1G8lDyUcN4BGu2i/WvG1PSkBPXte3LxPm9zTHJM3/H+kteWcJkLBBPNKVLdv0
jCmX7Xie7xKvdxf334fNmvBdS2hG0RSrQYSt1ibMKUbZ//9VbjfMiX561Jgwf4pQGbkmk18nOdRj
iSMDH83dcEsU09sbmAS7+WRYGWYXD2mB9IJrPEfRmwUI1zkAUfl5HMNKTjeLmMbi9POqF/l01HKM
gNr8zpSy1u1Oeml8U0G2w6kcrtcbHPLTTkDv9gyy8Th1XhwLWbiNzmIaQjBXfx7r0z0irEudeWNX
+jJ4z710W4FqX3PE1DjgaD42qEEBh7CGKPIaMghxmwXpnCxNIZqMuGv6ngfU6ts2PlVDSmn9fTog
FuEsPEaM44wC/BWng9VNeN87bXl1yK5ie8TngTnLbS6zIaJj05Cujb/2V/Qa3FxP2TM9UqkdQxdQ
e71boX/iUCpTdEgk3WbpB31SPJgEuuV3ooCqLpYvjrbeJZecKuRjNTIREtStk7xYXRXnMRYi/5ui
joyi4Od3pP8mzhkOtjwgSGD3SoH0EKbdYO+TnM6ciUVYEPUgv19sce6cgZJmsjXEh9m/e/h266nf
628UnIYiHHTPePzZb0QLTv8OfGSeToN4Kag4PUwaWKCzlResy9qSuhCgjJTfxeRmYi6IvNkNybJh
iitCQkK9ZAmaf/FUxCAK6kjM+9wRazDPfz7lfoMRuH6TTVUHG4aANIjKYM+wwCIgJS7s27mT2Gf8
gMQBLu782j/wGlmlDZzhJ7BpygaKXgELI+yDScjauC10xuqRs8sEBOt7QIjDhylO7bm/osTv913k
+X2hEZdPRdSyV/8YkfmYbtLR1hNNE3RAsRA9v9CYND3LMy3zkg1wmkK0kx1MlzNoHrXjFP9zDb0s
+daHDy5OxNv6/H6W7nl7J+odqan5sdxhVVrOTcxeON+BpgyQkW5SfbTFnBSxUlRTqISmcSEWkHx3
4KToV3fIqrxV1yv/xZiggPTkrCwZN4OHJexQPQG5HCyryruU9rEMUSjtCBJS3gPFtuw1pX+1LP1s
WpDNvjhu2LvwCFEGI6JCMq7ej0+vFhheeKOL+GSO0jN8UfqNQqBStpUHKLZDL4Bk+9hAcUxMh5uu
ZerVMIcG+YYfIeRN0bNtGtTRy2B1oriIM9F6z8crkKIO5wrXpkUpKLIuTJ90Xy9Tz/+S2YUhscIh
ac8ZLgKfAQSSkObybOtKBehPn5lJXbik7e2WqaeMwpbDl9BJsw6qfW+aLSQMu7TXRmS/UlcWvnh6
2eZ/KY9FGSrKHvrE3kW2SDIwVRo/rJ1GnO4+111kEQ6s5s0jKodKoczeNxKiMTQkqYB7Mf5+Nn7L
WVBj16jzvBfAM6n+U0iUGsb0Vq5eA6GYpx1rUGfQ3uOF5z/SxO54CqtyIUye9RpQ2e0qNYX90w7g
bT99SKhgwgf2m8FiFtRHI2+rwKfPsreBxhdDYgjGRmVpJ6WmyoG6bDyankt0dHsbCV8AsRkhD0dQ
JagtUgwkwsbADbnISs1UUKyUUjjQL905uTk+YNFgVr8PnCzvC05F2hLN6O6MiTDJWuzPFYc0EKff
8p133GiRZMij8VABTnchsdZQpV9DHqzhmGc2uFxrEriFbBcuY4nrcrc9gxPfs10DnZ8qe2dqxZwr
9DmGwfmrCgC2p7uNUymGQxwV7R+H2mT2DOhGXzyBivGX6/qfPF1GCA/h9FHl1vpK0Xmt+EpDP1xW
RnL4AqRhtJES6c1DiZ7eg6Kwua3aQyYKNrYf35qFav/D44JonpmvoF8Me52zmwR6rFXseJ4nYGOH
CEj9vvsBqFmxrUVOzd6TxdBMCmdpLptpJ0mR4oAqo6y+O0VN59oiPbIbjOkA9fNt6Alw2/4Rdqss
Hk3U+ZQb+V9XgvjhtwO4VnMmKwfh8kDtZeDhVcqZWEG0RZ8KmDICy8VSW54O7c1Nr84oZ8YkcEuV
bxfKSOUThgzVG/ZKIw7Z73Ozrfxtod4r/rO58zrnzCFP2MMMLRkcmbt/l/gUiDhhbVqturU65R5F
fb/1l9BDwZeGDc+PurZlI7Oa8tVWRzqMb9guyexVfRBCAMwVp6VlVuYY6iGcT6l6CCfHoo2vKk7z
MhMXv7hMz3UA3H00XdssAjEkmnncTcQTuOvdXiaSky5o6sTZKvalVzWjAuOV5TiRq3GiiT7tNRCD
vosIXeoyg0WbKP5BPevSNLgNZmfCvnCkGIRuBDJBvGT2NvBF1/KYmp8F64EQWANqQGIIetDGy19S
VlWkVL3ee03R+RIfIeae2SftuE68e3RKUWBYW6/n/Bv/njSveG3pzBOWeYOREWibViIGx05w53jp
oSEwTPkQUHKmYd68fpKr+IsfLBniQQ+guCHpzSXDzh7ry1rFz4updxqm8wUPgq7uKbDoG2Li8IXY
bEoGEi4xXw7N2a4sx4n77sLDuCjVAz+lAq543hjp27QGcmCJYFOVpeeQ5DOnme2NQ945xlD7cOOs
XX18E5UQDc246q1T6IAAoK5bhs1hKFs4K+kt9quxQVR9BonD++9HnTuY/bFIMeJEc7Qg7OBs4h3j
0Qa1wVjrewcEU6c76yBG4D7atd3UdPEhkCBDWMcDD47mgso2/pZQhl/ZnU49WHoOQ2pGH0KweeK2
GZ76VIgP5UERUt1aTjmvHmEbZSIYoIUbAoYPyNwyEe5wA/+KXXGW2J/VmOz455otxK1Qez5o3LkX
d+k8JeX0mahHpuoZuSnfAShJOHzzCVjywAy/a/kFdn+CCgBBoTE7Y5FNaOK/TWtru6WOi/WFVo/P
25LXh2y+xtG7ZyKtOx1MfMwAe9Ot1VkQ/daTugyCyQn82QhaVAYyFNg0B/wnt8/TTdZG3L6bcU+M
7EfSl7xjjczko7WAHWTVAPJJ+Tk6W1qk0j8gUnhL35iKU+3q1Zm/NUnpA8uy121UMYxGnVn1Tfud
Ui1CtWIT4vgm9wZrXYb9L/YunrrizAeLN2iLnFxe7Jkc1rPN0OJiytMsPdz4uERlwNacMnWMSP76
Xvf0yUbKGr2ntBd8mtEEpyHqdeFpbP9WpTGJ+RZYQeK2IlQn8X1is1zyhBQ6CCqKSeQlG0zhNr4n
9KpVE3u+Qbbcff48L3xypNH8ok+tgfTuS+F+MTUvIRhkVRpWhePjGq7cYPdRZdoDpEC3j6kgrHGR
LKzSONf6KtrHqvhD9OC2uAwMKTPrigNTxu9mTZa261zL2DLrBEOYrYR5ZC9rnnLEfaue8Sa8YkZl
M9zE/wwOxku3IjEgPm/P/mA557Dk4HXQ9QtwIJrLbAILmHGw5VZvRApBawrd9q8/sbbNIcrvDgqO
zxMnIyUhUk6d0zFI+FXSRQOCnI6hWwiULZUzbe/bitbz0oDMNwGg7HJbR1AlL7OtD/B7BOQcbYIE
yKDK2rnbU5vtSb2EJNqK4cnkv8M4uEVxxMZT2iQoPrWoxRUM6n58mff8CqlLzz/kgfkOBCMXa8IV
MTVTeYXuZsxrMc59Db4MNZG7tzACL2F0R+1D07HcHVfqohodJbRfqx8RD6KN3CPQgbYKejEqdfMH
Z+Wd8n+BZ501oZNGtZQo7SpUl4AvWo9YOhtwp1gTSo4aV+czNZ+1+/eri/SSYqxgbTO7n7VS2lOh
M2lwZa0J6nU5SOMkP+srF/WQwjU1L32ZJ1BzxQNwUdiXdFs42QpbWmKjfeARkkhFx2i8hzlO8yxT
UAjkn2vqnJAPkjxqPinR+kGzz2Dn/9F3N6IgnziULd452U7e9ZzB5ZsqrF0og2ZhTGpSKcl7Eody
70utVuXJcfjHU5rco9riLcvL62UkNJXMlodiE9cXkO68yUe3qzB0LQk2ff3a90GzUA8gFo7jCrpo
p9visPLStTHSMq5EH1dsvtK4fWp1aYyHRZktzhRC7bodT5fGBgUQtSWV5jDFHIt4mXSQzDCw6mm2
a0HFRSHTFmkQHMqAF/yPpe4A5dZ4QuZmYaPy4MiLuf9aaTd4mOUKc32HqDjiW5kSbsouMkLXduzh
Fhy/hhWaeDLTxKZLilsrYHaxvGdJffQHs65SiGV0acxcUTgxbaE5IARGUkFeqndhBvm56zDhk4uh
/E4WdKeh6dpzhPSBD6MHJb8SW17RS+hTqHavb9TBHddTUouCHKSkhIx6fGsvLysVFHV0kEuEMri2
xPpZP2oH/zGYWxt7ZJ+5ld/WF4PGnuU+yezWDORXjR3WuQADPQSsbfHKHADGv5k9IAjaLGkhk9fQ
GfLDt7cTi+d3H9yRHEPkfkT3lPYoIkhQr3rJTAxADWhvXBo0Cr7mQOuGe30qG0gfBuEmKPUNS9AY
hDUDh1CRtB+/ZjxTqV+LkiP1TudsrnHFLEwSCH/eiTvjv5K2lF0YQR+H1SyCYH830hpo9ei/oC9r
FkC0C0+qLJcLhz8Q/9imvqanhZRz8sGP9oGcYUAg9HlgXOVGxaYcn+wgshqwT9iF0kGXt8ywUl3P
bAyLqRJ7OKUa42Ohq4eIMDaBVzSxD2VJ1QrCGYdxHg6MUw3v6lFQCikDLnWGH+4BVd0SIgD0qim/
RxdID7JmnAAwKf9x6lKA7Vre82/380jmqY3feHVVKrYc+8l7erjpOYtdlskPCq4W11clXYnKGL+J
0LQgkvdIFdHx0MOsdiPnYSkt6w6oYvOYeE0fmhZBwO1ZLBuxBYoPcs1VJdI/ocDnx8VdDrVepjeS
20qtqN8fJfgfky8pvtftYhJ1xB2k1KpKkBcyJRR2tF+NT78ZpdYRSHaGu4q4WaolT7OwchS5MdWJ
E09RWoBW5kH0Cygue8j9rQbUoMNOv7/goMbN+N6NgP/ni0p0v/Nl/VypEikgJFg80FaySRzZpIUQ
V4EkR16LQEg5YZUL/cWzDmOU1YttecclKnVcGBlloe2h28FI31pHz2fPDP218RW8ero2/EhAc3hq
nk/WHYWoYdGqnJi1tHhuTU21pNX/azfGekHjFzXnb4f0rw9N7mfvi9NCURgMMadgfVKsRRVlKWjN
TdvikA47de5xHpgwvVGhk0dxadeYnFLvVp6xFQIkx479xpEXLCmj9NsxN5WA/tVTzz6aA5i2xjv4
CF9mbNNsMJIHZfyU2v6qcx9ETKw+R4IDBgos9CQZpDaGvWCyb52CRuFMnBBrqc4phg9Y4sPR2jtN
WZVd88ihgNTMQr1BfvD+UzQIH6DqTgMhZHJvm5VP4Zw3HjHRMcdkb31PKs2EPENbYPAgeSsLXJjz
MvxoMx8COuZMdK/AV94gsnd0ih4AntzAi7D1giC4U5INlQDmMDUJgsbBVJxvfBji9/Lw2/8mrlQi
WTwqskdPk+F4s2NcssWte/RS7ga/sinOTeFZT0QEPl5grFyjXPdtru1jguZw5gBDfb7hFKz4qrzh
I/waIDS3zafGjgs7TXcncX3JrseNIdtMLmzH6i2CApKPsfCtXuDTquq4Z/wxQEmmybd4ibhb1qZX
2qNaIHs2b5QxblmuMyX2FF8GAbnwcLbyCTZkOdief6/pX+/inaPWTTEZFPmL1oSTVkwtF+1OsMX/
XNpoqRD2doTs9mWRlGiuBk7nibRiUFTMOiRJbeAEH3SE1egTy5bx9C2eYkUSojHXCueHm3R23rMZ
HW3z7MXxkcHMRV4yxsGK0q2zcL46o2yMlaIArkI5e6tD1H5wJpUMN0R3KKX0u6/NXASoytD0ZgHs
2UsGekg0r6bA2aI8mUudazqbYHGZdEbkOVIx98Lhbfr7Z4YlI1Bj9S2f5t2D7j+AahKyS4HeQIeH
q1guOCTv1D1pqMDiRmTj8PmFKiUp3AesYtwxlroYDbz6wz0TFQUpr10UKB/SoBiZlN3ftmgAgb3U
A+BIORYRYL6UBMpmYL19+lNOtHto2XcPV4OGaSMINcXXoOJh69ZvHTPaUscm667+AeW5voZGXV4A
ttxjHm0e6grWx5jlhWfehZWNck9MzYeT9OsaDO8T8YiCsuyqshqwAEfFfzuRsJhS5+pgAaiab1Ef
I5cKW7GMJjYeGtMPavGCX3ByTXNlbDssQBqOb14eLdXglcqqTT7VehQR37WuEvGRmsAgWazLQmcF
nAbMpAb3mGLHldTIm2ZGFt1WbNhkVz8Jej+GTurFt5oG9OoVokLXlrNfmvjyDELbwvjw7fnKomdg
2tAEZp3Gzzm1bL0QhLqnoyA52lbf5JiQKcFsI3rcnniADKMYudBV6w7JQh6jcBra6MwWHm7yQX8z
kbxPLb8qIllN2UB96+HUw2JJUjF5h0vQ6wOdEjjPI7ECdI6O1qG/y8u7/AGa+xGa9/lIHbg1EZpL
O6NqXtBP4DWtAhrspx25fZ9dY936LcEUD5wXQJzeR58WzrZVWkZflw2qwym2Rzdq6Y8uQMGLdUI5
o0GxeIbCj2UDxOIv3jKaKVVohJQveu9rUEXgOORHGAsECIS+qQTvcWFTIbrdEU1lOGz+644kOHVN
knTwbJjT8O9+i1aaYFgOm8N/0TgHpslsbXKme7Yo0UJFxeXUlJbCkCaTjsc1U3wxwuhVp0U7hScE
V/H2eUvQxpi5q3bFcs6APRHujarusbffD4vnj6TlOst7CS9h7MitCRjTZLAnUJ2J4OddM8W10Z10
KEVCFHRF0puL9SVX47o2/d3eUJ3ohtYxssH2EvdzN6szToI/uQLGbbuXz5RXOnpMQF6Kex5aLYCc
9IKasuU2ToJ4O0TyXF2vXBuU1eZgujPBPfYwkqFaG0kImDsZt5tu4s97fX368M61wasfCxwkBDUb
0jLByGRyRL+iy6XT3mUOilMy1F+qIKrovh0Gpfs2t+P2zCl5tLOX6RBr2VutGYfve/dUEF2T0xXL
Fw9RpaCuSssV7PDAwkjskC5C467I76UmPMBhUWzJCtwafgymkjJfS2Q0+QTomHDpdofmEHQhMXij
RuMhJtzOkJiY6ZqhfpVbtLmEZDsa7ohwAI0ohNdAf1malKsO1d42K9n6pOkzWighuRFmBTgah2Sg
EaQ6lkN+jrtGDghCAotiNM86xTNNd4UJ5DMgndlZTxUds73uaiLmj+OWHnewQoC/1pwMNAedeQ74
c+QXle5m+yzxghlApDYyRFgxvsHWnlzxpEYlZ+FvD0/jnv5JZT5mqleRHtb7UchtN14f1zKb7rlm
+ruc1L2wTPzK2ZTHEn3H04xOTx5GjeBQed+TXdj/YhaRWbOgmfwDjn085GlooL40OfA01vZfPGpy
/rBOcMgVGAkv6lYGOH107dd/Gzk9sQfNUEXRdxYOh4poJ243XENpg/r/AiNjpPPhNOabt+NW6P3B
2f/wMxnHfOmad+fcn5qet4eQwpjLOXxTbqPIvFEfQlpevFv/aA5F6GzA0y1Na3BMp4QA8tQ2Rp2a
DgX4LJzhXgmpw5QYhNqy6KwnDwH7pLuTCJT74zvrKjQWZyupCdDvuKWLWA2tboawCdDRmkRTmBGt
YKg0yP/8z9TSHIv0w901TaXdJ6kfOOPV2E+/NFJUJEB3WfJLpucNdsGmsK4FyAxes+mR1KGQ71yh
Sn6YcX02HpXVFD+1m2xH7ICUwGTaVfU8qlQkm24a6Nk/Y9SUEn3ex6ZRebpF52BNAr0IxojiwhoC
tD+IRLLWqpg5MKZNLiZh3WTvyIuIVSIGVHwqxoI93Gyl8OiTuPjeTH6bJ3oDygb2XI1ws+aQAhzS
vDD9lEO2HONUYA5f8r53dyYT7jdiNhNXt0M9LXOMQ8YVSnKLy+302iaNYZLAKPolgnYdPughE+GQ
ZeCxzAq3Agkbw0xwIfDnz1RU3E6T1GSL0xa3k/lty8wUVAnzJZOOsSiLwe0zy5KywZPBbuiPpmsK
JavmNmrsgOS6Z7GJS0HM64oXWcu4jT1FtIuvRihsI/G9FCGPBpfeiQPkJngkRS0Cy8yXwRrVBZ9W
JWuU4ZN+5Aj5taVedP3n6AvY3l+ITTbfmPFJdu1c8A5MlnlYZNJsVw/qLFIWlB2DZikIJIj4Eefy
BsW8um+jR5uzcZLr/jlSRyHWdCHeHtciP3P8DxDVRxWmqdiZ7/ti8PBpRdb3SqZrDol8iOoDRsA9
DdKzEMp13L29F+qfe3j8vbWXFMAM2EJmgZdr6AvNVe2Zw0OO7W5TMrwER30AsbRBPnqYpzRd2fyl
JMkUrNOoZOoygKaZqmbKA+OjZUgyhiI5R8JT/7QQNxT+Nu9tyPjSjFXlVmU2B4WUjpQrbDT748Ri
PqXI7BtgYj/0X6dG4abnroKIR8leSKaSi6wWtkE3aE8gSZQQUuq5tUQvR/gsSXCvvfj09VlatQoG
2noHCeXHHtNcVsD/i4B91pTK8p+4kdEtmPRXIPbpLLrhOOMl6FdCc1RuxoYSFVS+hHz8ZHWI2oUu
3PZDyRw3cT8qWO+j76lBuDEfKyai+e1yEAj35gcM7T7/uKEO/zCRDCx1cVjNTafQLJF93RI5xWfY
LzXQQwtNAthklNLLfMDcruGc4ClcNAVulB2peOSUY3R6Z+nPo4WeNmYnIrPIwCNPzKp9UZWNA882
QiOdxapbeOth7kxK7RSgvn986uBlMpknBYmET4iFuoFIsQwLN4dQPSGW8pOwQBfN9UQsFx3e0qbx
aic92y7eocFkLO48VExQRlOvtoT/OKBk4wUh2GFMHor+TA7XlPPZoLV3Bzcr3DGAQ1SxvwC++tQX
YybSvf1TeCW4FDv416f5sM+bbGHGIRB9EmDRjou5kdQ4/1VNuGpO34hHNOmfJiPo/4w3SinePL4Z
KuzGmrRCKyjNR3PaPV4JQx76+IpZraAu3Ydky5gDtUNsmzmmq61GZfHvd9pwurz0nkuugJ9sroi4
3aSD0wqlS9G5MFMf30nzb+KJp5Zvf75vr+yrMSjNNxSnQTkE1fv+GfMRRlJ4+60tpVO0HvRyVsLX
bc8TuOYy2lW1p+BqBjKr86L3QvponAMeHdTlsXrnl04G3o1bDQ12VeJAS3Io8Q6kRnhI11ZTQJa/
pUL66wwQIiXBziuC5uuLoBsTAr/r719utodE4LinVGyje9BtqUncFis4FmUu5YUs+DirN8Kpkg6c
Qwdinp9cewvXbKRIKM3IVmORaBGg4NePx1LcLmyu7yHiXQH/SPszsVkNQLFF+SUkrU6lWV9Qp64P
fEuqW5UAOmGWO2DX6UP5EmuPvCcvDKCgutAPfdy2aqqq73y/MR/1I8unsx63LRyxJWvRfah5B8Pg
mt0IgIXPzJ7cOky4SFWXoTVF+qzmzp4DtQY2bbxUlm92A7dWTZgngzPS39Q6TZIuatBVHS35LIHi
6bdOpQT0PeClYl0Yykiybd4DmRVylRRpx5CLrUEkYdpsuKSFYoPQyBJ/nyJrwINB4g7kYHgmaPwJ
6f3iSzt1Mo3WyJMALPnRHFJU8FX2cGRpK6pGpBxsL2Z8DKWQgbDgxH0h9ueq2SxgD9zhBldSqhn0
l8+PSxVMqcuNLoz3rVd3Wi7mAzomi/8LOy+LWWcKP/kleSmDDCm0bwShhgubWh0pV/i89NQLYft3
7aBZId+eVwyn7jKeH/OYkkrGM9VU3QiB6n+JIwqIxd4pyieJWPS6VqokA9xv53VmZj+VXWrcrj6C
vOGjaX5sTWm1HPMyp8mX9z+zx08M5o0QoaaqNQqzLa5NgtfAwhzR5l5G15ygNzwz6dluny6oklWG
7fEBn5wROMJCcjQ3eEgPr2mm7O0mO5KARfmii6Hh41rFJogq9xpZRxIb9ZIGHI8DcUbbovDdLB3A
7FEK32iaa3/rZ0cAf6QxRjfxwnOj0WemM/h9QFttw1ITXCXJF1OV5JdJ88w5fQC+eszE++CfCsCm
tx6izXYVn5J8JYA3GEMwv8JR/QPBkP0CHYE9OxiHWdNdsz1/rIn/toDd5iJcgR2LlC/9LExkOEQV
xYcKQRHq/VSE7Ul9jWqHP3a6IQcK1xHX6eSFUkpmyx+aNRhzOFMJLIczeHI3+0abqfFwKVswO9P0
IcDk3Q7/TMp159kbcUpFsd7AB3xlwEa1y9TN9fvamz0S7DG4LDmJjlEmnAY5Qax5YoaZo6LuwWKU
BJb03WjUZTsMnKV3zBBB98DgBxqlxjSIEp1bDvPXObIVDFTm0r6yZ3jSyAS27blCUbD7ETkAZMkx
O2nSla7cYC9603xbfwrYCQNh1BiwdljxMG99a+r7CQNCoG/Vt9JaB+ku3qFgr+JqzKLWEBAVHLgU
hTj829Jqbo+JPcV/RxTU4j1W8uU3mgCZ13hrHfruJ0epVXe/UrSeyC5iNdjSy3abTpnpdmZTo+yE
/aHAlY97I39Ea/0UbNoB9AiOPYvYmUfiXwpkA3+ngbs1hgZqQWyAtwurSOMrHbyYe1j+I+QXjIJx
WP+WJsb67s/5Tdv4mx27q6raDLsP2S2TzVrvayvAl/plmSUAXQVI74+hCDmA/rH+kk0IUpEkD2nR
1sbJURj65qaIRQGfNwYaQRnJkuS7eNU9k7tVhbys7z/5YQ==
`protect end_protected
