��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���l��o[��ɴ����>�$��	6������b@�	������b��VJ�o.y����L4���Z��1룠������	�<�~���E`��-�R`��k��-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_d
�t!���N�S��گ/�TNM{�C�5���M��;����L�S�:�{���\p<��)�0W��B�R<Qt��Ԁj,3Ӂ�v��`s�HW��眣�U�Z.͓k����W�z�N��VXi^�p�ޒ�}۳ù3���V����U�,����[�M����6؈�О�X�.�, �|T)�v����S�����.f{��4���!+t%a%U�f����b��0����.��i�tn)�Wg����I���X����O���� ���z.�^q$Rc'z}~��%7�~��s�A&�"���R�uV<��8U7�I�9$^�pz�w���6%��i�ʅ�?}csw�ci��ӟ�NA�q+ob��{~ףM�"Κ��m~��T��@�VRQL�`U$�tS%�m!���q1�(�"�X�����O�Z����~��Q�2��Ó{ �WB�R��q�|����Q:{��:e�ϒ*��ahj!v�~ �4.4W�;����hOp�����v|p��!�/���[}���]�Mq���qm2�_��>g���n�0Z$�μ{R������̭l����X<Sd�O�doX��΢K �Տ�Q���ooD��>�I�X�˸�n%�y6�3*Z�6��B�X�:�����CX���`�������(�$F��:�ܟ(_�"����[�ş�,�y�@�בּ�mX��~Ԥ^�L���K�^��0�
a�~R���.��J�!��ڷ�-{쬸L�@����}k��y/j�K*C��6��d��p�K�C)Z�Ƃ�݆c`K�Bݲo��Bgp� �D��	��E?��ޙ��|�7�"|֘�JR��m�QY��$47���}�k��l�
k .��������q��g*"u��A�_�3ּ�ʿL�}��ű��l.31��D�Q��c��l*f8 ��k�X�d����j�}�qO���;��u]/�e��}hD�1/��!�$�;H��e?����|YA�(iSOu��;���,J�GcA�<�<�����h"���������H����������}��q�/Wl�G-u���5�����I,v��/�[5��OK��;�Rb�ȁ1���:	lƄ�-1+��H��y�ȹ��!#~�<�,�A3Lrn���v��&<�W]�/�&���Z�c���������6�`����c�_� L���t��!�6���}eѨ {���oӁ�~U����Jx4�l�Ķz� ﳜE0B)�2��͔Pan��U���f�ZD����scX�h�T���V���ur���@~ε:��kV��l�c>a�Bk�g��7>���<@�y읣[̱1טw*�47�|�)n��э؂�.Gg���)}Akp� �!�Ew=��'ww4�
���ls"��t����E=�M��y�+����7�p�=��_��1m�	��27t831a1`��e?cP�P.�2}ָ^���?k���/��S���8�U^�Ս����Dܢ$��K���wF�gd�ƣ*��a����ک[V>7L����+��lp��5o�y޺��0�֡�'q�m\;�y����j��n2�&?��6��h|��A���u�9�P�X땾�����C=�g`��k��cA��=eڻ!�g��.�#����\���7s+�����GB�u�tȸz��e�DV���4�B�bKVD6�����XcۢDpŖ�"�l'�FV��`�4����_# ���zȣ�DF��:�xr�+�uF�>
��ߎ&�4��)���ם|;���M��Y��L�`Kn�^?�؊�r%!9e��	I��ozt��O$E��ٞ(��σ������<��B��O}W���]�1Y�l0 Y�῿c'"r�>�� JJɘ�\����RoDmw�-�u�<���c�m�DR��#���C����^ua�qS2�ؔ�y�q�3?�?������C�D7�X^�a�2c��B7oɅbb������oY�8�Q��²�x9�yx��]�dvc\�?�%>�Z:���=��g�jޑR��0���M�������.w�-pB���k8�o���t����\m�m)�O�l��1���c�9$��$S�h�� �T�͙ 	� Ië�����c/���w����E�Vy:u΅w9�1r�j���?�p�
�`����f�:�����7v�%�R<ve����d�C�@o�pgD�Hڸ�/}�D�Su3�M
H���A�ޛi	j�w�,�T�����e�{&1�V�4��L\	�Ж$���?��k�������hqu�?�Vn���ӎ;�6<*S�v�]:TĘWL���x�	��B�0L���Y�n]0j�?�����4m`w��cő�0#9&Xկ�P�}>OZ���>���<�	ZJ���/K�q=i#���n�J4�de��}���@�->֯w�\�.*E��2��T]Xo�v3h7��&�Lo)76v�$Tl������b��7\tһ�$�b�ԗ@���U���y��)��Н^ϩ�o���}z���{pa��������
i���#?iPC�~��2���Y�?v"���v:gt�`�5�A�+h?d�*��շT1Gt��������
DS5Kh�W��x��x�2�/���¤����d��h��`�D�ڦ8�Sn�"˃�x�s ��+���ޙU�:C@�\@7����4:V�Ɨ^D ԕ�φ@�"��t�n��O&1�V�mDC��Y�0c�c��N�74��>���I��.���8�Dd�?�"deW���ћ���l�.z+İ��U-a�lꅢ������64|�*�Y/�����������i��x�'3ؾ<�Q�2iЋ �c�Bs����l������x���?3�������D���I�'Ô�.Vu줘6�7�4��Yb4�h>���Q%� �}���W՚/)#E��_����ǽ�} �)����zwW;���%K3�4и|�0M��O���^�-E��<���j3	�-V�وP�0�����(��q3%尦�>��+��!�F<�K��m�b��G 5a=���7���P]�� ��7:��n�3�����gI�x�Ow>R̚,�E�^/j���>�WO��{�hWo����28���p��1��	y�y���&XY�����O�si*]�p���vGA�+���".:pB�-�W는��\F1 �45�3�(�&#��t(�����ض�Y�j@>$��&�loэ��x\߇T���aK}\�uʗU�J ���C��45u�((*��>\bp�s�P�+x���c�
��L�A�!�	iMD��, ���("��op��=�����������ٸpV@N��X%�`��0�*:h��,��Vh���g�T6�|�ěm/����U}��T{��г�B��t�{����%�����h�V�s�ַ�	��+/�w��AlP�.7
���šgm��L$���|�J��t��ۆ�Ͷ.l�;=��m�D�따����ti�s_���{�;���a�P�o㭥�9$��jv�Gbތ�C8��	j9/��&Vp9=S+�������ْ�o�=�$9ʊ�������;I �U"o��x|ԫ�di�|�N�����G���1��z2��*�I�j,�,���l܎�9�W�D����|�A����ª��pPf+����[c�uy��!A��+n�,���KgM�P;/ƋI��t���&� Q$��|�Y�u����a�$�X�^��nr��}�B�GDw4 2�������+q��A�!�-D���nN���Ņ���Ft��`$Oj*rN���6/�;�J��*��L�8m.�����ǡ�!��`t�u	���4���
ߛ�T'[&#n������2L� m�g߳�}�T�����mi�@��u�:���@Sz[��>����rŠ�4�4�G�. �M@KR��u/e���I��'��Qo);�n(v�H$&����F��Β��n���k�	�\�z֒(w�e�s��	���9j�U=���Y��ݞK�}�����E�2݅����Q�b"��F�-���%���I��[Ǥ�����%�3Vb��kձ��ҫ�'O����c�Hn�S>�~�u��E]7��n��c��`�R��d.wV�L$-m%ǩ��9O�%N��'�O����|36?�	�1� �
�b����A�|���u�dk7�2�A#ؘ�z��-w�d7����%-�;GA�� ��\D�?qڽh�X�����8(	����I��{R�6Ss{����#�ι�/���_�3�g��߻!+��+	�oL*I`���ee���; ��y��} d'T+c�)|C�3uL͑���3�@�*�	�����!n����t^\��
R����$�<�q���єۺ�/�삐��zʓ���lqF�虤)�R�� �C�\V�dP!y���� �������R�U௯��j������KmD�S�}�D�}�$�7���8,A`�� �v6l\��v� @�B
hӕp
b�*b�z����ڮ�H_�%�K' U���OnF��|��g^�+f��i�VW゛����'���y��B�Q߄��a>��j����Z[�*�K-��`��h�u�v�wH�b���~�)����ͣ��ҵ)Ų�C��Bk�z�iO5�{��O.KEIy�ځ��Ɣh�P������+��G2�@u�9�����#8��y�����s_̈ѥ%SSE�A}�+g�!����L�r�Ax�cɰ�u����x�_[�w�v(z�@Y$���;|vQ0�h��QKk���ڲQ��R��i�n�����%��}��r[S#�I)��»��e��/+$D_%�ts��+7��P�`��rK�)�3%��E�	��6�}��g�5�5�%���>
o�x�{>9��{I�$�U�[~�����vX+�_9>�l���@��1�L����dX�T�7f,�;P��X���`-_��7��� |�F�_��QX�&�sX��}ZbA��f�H�NGJf���;v�WL�Y�������b��P]����/��:��m ����'K<~��{$X�D���C ���7���9��ٟWF��A��dYT�nN�|�V���-WLV��َp�H�����R5sօ�yn���fǕ+��l	h#��o'�g�}���`� ���b��J~�{�K��4��k�=�a��1_t��}|��E���@���a�����k��10%�ׁpu.�-?�N��e������WLO	U����kɡ�������|m���>^Q?�k; OK�C��E��C���F�u��M��ȕ��@���xOd*���tU'�Ý��etu[����\��W���P,GA�}���%��o&����:�w��1�`JJ�O!�d�g�	5�Y���/��0B=������X�-�� ܰS��\ky��J5���-�z���5I\~�r�x4�}�Ҫ�A����̲��&<^9�^ZN�������x��1Y�+�,U�v6�˶Ь�Ĕ
������i�����c�v�J�ΫZ���˥8c��C�89Õ=2n5�e/U�)�upWғ�|����5�r�jG�a�Ǆ�hB�l��p)���÷��M�6>dDy���s~��cg3�sv[ѺC��v�w��w`|K�=G�V�Đ�I�BX9�zx�1X���w�6WU7�&�u���Q:�}Oct��/N�Qcy�-�����-(T�"��_�s'�LN$���^�p+��s�r�SX��BPp^�~5�@Аc�d-�ٲ�9��wiqg�j�N�gf(��6�ՋT�5V�+���Cf`�j���
E�An*����4%���K�N���>�R�FόK�h1�W�4{��+?�x/)'@����Q�+�ꣿ�;q�H8��&���\���Y%h��(K(v�	�R>���1�s.���d�0������� ����$���S�r��6vE�Q����31o�Hp0�����A�O	��c5(������|\�x���\֎y������O7QD�4�qw9��b/���'$�&��b
�ܠ[#㢤-���4 	hl�n����H< ��3`mu�LZWפڼe9u97ݧg^>��|�BҽpZ�_E<=��	��wz����&z� ����ϼ#��-����l�9wʈfn0���b�&9�� 9�[qskI<n|��qE�H���ʗp���,��;�Ǆ�}��S&]�#x��H�ҭ��x|�A�t�-�(�KH���)�b�3�a���c:م��y\i����֏��
#����:���΄z.낪��A�;�WlM��"�$1	M���I)'l��2;i�L�A�ź}l��;�Zj�E�. V�Cy@B]0)��)EԜ�w{�[E��z�A�2�A�w��е�D���Z(�Ӵ�
�s��j���Zk�RY�D�0U���S�T\��e��JG���!�4�(Џ#'7^���h@�B	V&�C����[��_��������A�A��Dq,�nS �l���=�@SCs|�z\��S��2��6!x�0[�O��8���k��C"{��U�Oa��vƿg���r�ѷW����i�����L�kDBQ�U��� ��:�":��GJuwB�]`���ݡ��H�6���Gn@��|�Yyj�~*Cd���
�X���T�PF�0{y�����ۡ����j*�ڵ��X|�0����8ǰ����z�L�t �[����k5=翇&���6N�h�g�=���f�ʾ=��~���`j8�n�	��V� L]Y�7�Bt��"%E��E��鱊�S
ƙ���zՕ���
�m�*C���"LD��_�Ќ�?v�!�_2?�y�ډ3�����[k�suX�.A1 wH��Kbk����+:��P�SS�o��M�8��dq+�,��ãR����S�ӵ�@�k�w��G�����@�4���Ĳ4s�ugK 0��V����A�~Ĥ'���]ͺp�	;��Vl1%�'��R���'�;Yb�I̹�`g��Vy����"��uV
���Oᯰ���D&t�Đn��_l������Z݁�����ޮ�I_Z9_b�l=�l�"����x�r�� RZ�pE��kxo��:�{�-�+���$��T(x���r4Z�Gq�!��0���̯���F|��~�[ K&{��3��"����z�P����N��'�2U{o���Q����b
�uᴲ׾n��e�/��$Ƿ�ܗD^� ]J#���W�B�,�����\��Ro�yu��ݹ[w�:� �7iEU˶�LңUN�ZO@��Id�6j���
��cuؼ��?���}�����gk�3���LЋ�d%imyWG�J�k�Q,C�yO����W�o�W`b��d���R�n�Jv�[�&_�����aW��6=�����D���U^6y�yRV(*q�W�I���=��t��h% �26,���a���Ryk������,��qS_�a�R��G���$����DV ��̘p�𔂰7�[�'���NW���di5�ӣv��}�����Jyi^�g<r`�	������i
L��q�T���������:�.S���P��y��+ί����f=b^������U���ӭޕ-��G2�?-°�G#T����Py%�K�����	凫ܐ^��3	Dco���� R�n��s�b`��#eEQ��` �/�4��0u2��1�7B�k��~��;�.�����g�dH��gp�(
m��:�Rnh���S<��M[ASu��fmG�Ѷ�~y�j{o��	�EP^���K}��]���&�н6�\��uW��Q�M��/��c�l5

3����=���i�� �%����
����X�	��1���h��?�.Iu��{G���>Z2�$�R�nS�����E���'^�{	�M��=|J�:����"��(0 lT�ͭ��b���/��%8<���7߂��lN�8h��$�V�H�#8�0�����e+�I��������6�	�&$���rϋ���EAy[�ҚV�B%@bd~���\����Gmn��l�ܧ��Y��c�5���g,7sim	6�����BVv%�
��0�V{��+5o�n-�Ӣ�|�!��y\y�������|�%�R���g����x��B�P5Ia��q�a���� �:�F�����M�	��D�@���I��M��V�W�)S!`��Z�qQ�0��� �<�b�	�*8��Y�L�X�� |����eow`�DF1���
���c�i��2˗o	:����Ko2�Vm��d
����}�@�Ѷ�T�-v$)%���������uH?1�g�.7
���I#�,�b�3���I�׌�����xwf�͋$����|MO��7�"ή�E��XF����2k�������esiQc��r���ο��)�;1ۦp�,���s���� k�{��#�+� \Qt�m��YrBy��(�oZ������ �-�i�>���a�=��h��$�����"/W�Y��b��Q�A�o�K���-
�-�������|������ǀV?L�)����"���T0���b���CE�luR��C��փ�?\�c�q]ꅛ��o���iB���\��\7x��v��@����Q��kʱ��R��@�>�e	M����t}�3�Ɂ��"{Y����lr�_�m�����Y-<QF��Z�@U�<�����ZN4��^iP�c�:`K�q�&W$s\�[a�NpZ�X<���=��'Ո�y��:@|a��"\����Ե��Ľ�":L8������(���z���
���5�KM��Lu���_�ǰ:�
=Wl��K����o�� �V�>5�~���)�ݰ5�!�<w�c�l6x����.��=B{�B�E�[���T	���HP�"F���i�sz���g���M���E�k������7�&�Ǧ�]��t�ۮ Ýz���仟�3@���=�[�H��e!v���L��-b�%}��P��Sd灮���}���	���Q��f팿�
�� ��-)9$jG��5Աi���u�{CZ2 Y�u�G[&OVV�8ȑ�c�O�#��J��*�փO�A��n!l�`�� EX,B��S�T����V6�W.#�W�g�ɾ�Ș �{��"d���m���*������������ʊ���E�5��L6��S'������H��2�@��Q� ��L����x�<���y��:UX�:^�s�Ӹ�'���]q�MG������kM�U-�nu,b��5�4l	-����A�����S�F���\���������c�Ժ�A8�������)�9����i�\�+�E&�C=>�n4���Zc���ڻ�^{C�Р?���!���0aA��T| g̼�'�}�@��,RQL[����>w�.v��!e�kԏ�qg�Q3�����&^����o<Dm�f4a �w�8��rƺp���z����v�q>:ui6/0�B8v�_�az���%��!��1� vz�yg�Z�OBg�[��N;�1���Gc��y�MM@۰�O���k[=u�Wd-�o���P���{��m���ME4?!�[�Z�7�[�H֍0;c���?ԝ�3Si+��8؋��FqZ���<r~������Ůn����B%mދ�K�%%�s480LW�ы`�E�P$�:�eޡ��5��E�9�;7I�+@�P$Q<Zgܟ�2K�9y$j={c�n>�����'v}5b�n�E4��&E��>�y5��w5pl��'̗857NV4b��P���BSb
���`��~_�#�D�-p��Z#]ʚ����8����'�����q�5`��Å���'������\�q�|�P�8ST��y��m�e0�~I�y���>g���Ս��X�e2Z��7SEr�G�^�������ݧ+�U���Q��xK/ƀ��>���ad����I�z�f<�� S����ɬ���C�v��"���D�EHxOvj�i�b�w��bFS$�m���9��f��1�	��m(�6{�ؔ���c����������n��v$pl���.�<�@��&�;�޻�gb�wd�� �淨(#��G~.���Ș��X[�87�ӳ,�{�Wu!�u��e�fN9D{9�����I�	&#�:�>��29晣Bwb�D
�"��g5t�}�rᦒ���HƂbR��0�Of�l?�j����{�yK*=]k��y�6$��ϳ��38�᱉J��PV{Eyl��Hh
�^�2��-Nh��Ho�4���;�fэp�	�d?��t�ዡpA-�غHZ�_<��i�w]�OHz��%�c����O��X�C6�$x����f��5�a���^�.�:c�;]����6�Y$1�;�i������&׀K�Z��
��qb$֒*�--_�ɨcsO����&D�0���A�H;��\HRVy'��	�U�t\x��Q��r�����+����8`��|/u�[W�?R���kS��i ��װy�t�~׵#�����$�́��(i��C^(w_^��{B=%1�A�Ԙ^�O���C����i}ۈas��u�7�퀅Js@��R�,���a3���8%���$��Я����U@�OJ��}2v��T΢C.��	���+�L$MWD#fr�*���C5���K�,0�O�n���gg�F�h���</UP������u%�ߢ\w�cًl�s0.����j�|�{K��J������Q�]��C�O�e��ԋ��+*���>�2�	g9�W+�m�m�YF��e��Cj�:�3{Y���؜;���w����%��f���E_�Wrk�z��E� �/S�0�d�]��֟(ܮ�h���[����v�iK�f��2��5��}^�r�������Ew�M=�(V�ca�x���n.Y`M�wi�SiҬ���,�~_��ɗl��o�Ժ컒��7�*���o�2��Z�~�4h��|�۾�<��f�9<|kdVX��?M|Mv=q_f����rGZ�y"+z��k�2.�ȹ���N�pOߴDX��H�±@����Rs6� �y|�Ll	Q@Af"لz�c^6����DBc����/״'�JS����X���P�h�K��h�u����4��7���o��	��4V��
�o�Z�!͓1ë�\J���|��j�͡���&"S�j��3���Mx�V��.�)R٬Fd(��r��2�{��q,�	���(]1/��'�6��w��z��Ǹ ����R���b��<��&�T���p����nM,ͽ��oR���MAS�d��TF���!�|�ģI̷�*'�~D1_�=s������6�	g[�Mb҄a�u*���Gr��ub���F	�w��a��76FY�E�:����Tc��'�'�*$ck�/�a��/Ѵ�+D���֣�d_G�صi �U� ��jT���}FS��B����6Jw��C}.�B�o��o'u˯ې�Jq�~�}`��-�>Q�x�k�=�W6��WӕU;��/Ikl�C _�J��� ���O�tVmS��g�a�H)�3�liufr�dR,�?ez�op���r�M��ߞs�;��r�/�a�^J�N�s�&�w�#߹��{��l-g�韛�� b&�X"���b�t�[k�:K�M�@"�
ce�� �8� uh���+�q[�DFz�'���k�U��B��+o�n���4�g]�סZP�������-��<�ޫĨ��3���O��D��K����J��u���
ܘF�P<n ��9Y��\����˽�J�7�?:�����[aoM5*a�)�D����8G��(�&�fR������4wk�n�p�!�o2f��j��ֱz0>&��E8[�{(/-�� ���;�.���˳Z9���eA�Џ,�@<�~g�G؎`�E�r Q2��]Z��9�!jΈmO{vtԕГ��01XaT�.}~ͳh�T*D�*^���ד8Sa:�" ��ω�Q��ʪaCG�j?��Ǘ\N��v���]5�P�L�;kB��-��1����\`	�w�g���"S��w�c!@�� �3#���"㐬k�y0��ܳ�~5zj$�?�����d�og���9=lIl셷,K�%���v���e	����������h�ǿ0���N�.�f�l�%R�Ą�eJ�YZ13j-����t��9��L����m-/�ˍ�W����y�TES�2fK�Ks>h�k��H-�`s�#�]YԿ<Ԏj<p`Op��a�l�Ҁ�����mԖ1��}�g��� %�V��L44j����hl��l.�Z*Q�O��U�Mײ�.��f|�:]g��h���ω�h�b�| [�rCs����d@���mr����e�(=0���~�,��:z��OB���e����ft2�5��d�#ǹ+G��k�K��Og�,�T�n�ϱ[�ȸ4
HՎYKB^�{�ʎU%����7t�%jx���T0���ͩ^�7k�'<4a��QS�?��϶�P_N�R;�{bD��o�r5q�ky�E����=v�����EZ�����4Ӣ!k�WCK`R�O:�L'H	� +�l3�]P|�yl��B�v_I;��T����΂������M]	�z+��U����E��'Ϙ0b&�؀4ɟ��k����Gx�\���5���d��Ï�tV�r:XfF��W~�#I��Y�gjK�eGu�P��D��e
��ɡnwl���R�ϯTF.�����h��l�f���ma��?�	CCP7m?����'V��g)E �o? ���I��DL~e2�xdg�Dɿ����� �e��Fy��f���_ s:�XY+k��T1�TAh��9����I�yv�qw�`*�)���V�	8��]�l�ƚ_���\��db��r�9��F gX�B�B��<��n1G��!����Fy�CDS�K�9z(	��F���k*�ao���O�<M��$�Ѩ�5 ���xv�2b2�R�9�~1m}۬�zm˙�.��c`0]f�w�j9�K
ml��F���s����}��{7��
�CT�>�&�_J���h�b���.yP
��s��c	t�����u\������xev����O��tg��z�쵟`f|'oN���2�VBx�98cb��+W'����M��#ii���C3F{��6�����$s�]�W��+���T4� �Q>ل�w46�S���ݮᨄ-�3
�}�F�?WD��D.Zy�ϋ��+����2��A��o� �#7�4+�E�4�ܙ<;�l���Wg��u4���e>!a�L�ح:*R��
�L�喫��0=%[>��3F�dn�_j�=���Q?��Nx�����F��K4\��v �j7��f?F2��R��NW H��%����>�۪�p1�s��|J�QS�œч�ؔo����y[��!4Pgmy��NEox|�jy	�IQ˙W�zw>���ں��d!Q8�T���������h���;uH�Y�>����Ը���9��������̒-��K�(Cx�G�}���W�-2�Mu�@m��xq`��ͅڊ�z���#�iS�'�ω7ؔ�dK���,�Ka��tp�<� R>�Ͽɴ���enT�셄01Iu���"��̍0��J�g;�v������ƅ�ʌɘ.'
5^��l��cGھ���;L��`�/B=��=�)�	�u�]_5�+�:��~,!=�|�����Fh-;�!�b��J?iX�L�Ǥ�rd��&}��HjluH;X����q����>X�2�P������0Q�~}�P���f��w�Q�@SV����	S���F�k�t#B�C-���f�����ɳ���J��/��NCFp?��}�.V�L?e���-s�A6Ι ��S	�%'"l�`J)3���k�'9Y��^?J�n��,n؂ώ�\��6^���������1�\�#Mx�9�}!���D.����m�'H��a"	Du��)��7��,�hM�D���(��Ī���dpl�>��)C��L˱�r����r�c8n#M^/�[�M΂�z���P'��l�͢?5=Yc"W��;�dT@Cݡ�R�p���]hp�Ҧ��}:��Zy��C�ŏG��A��x��wVߜz��4��9:��{p;ܹ؈1��}mk%�0����c!Tw=�s���1���!� ҡܣﺕz>y��u�����_D"`�hq��@|�LHؠ�&��euQ�U$c���V?��*b4�6�vMd�S*Q�|^Y��GPF�T"]��0�I��[W�l���#N��TM��ݲ�'�h`�N*�4p�2w��=�5�b)�ҹ�p|�ԑ&��2b$DƂ�Ħ���1�O��f��ArD�(!8��A5T�WݫD�y&�2#�mQ����PW�4���� y��g%;9pG�7���lO{�#z?����KB�ZW�F�����l-��J)t
��v>��zJq��ݼ��UfP�&��3��8�\�q�:����)�*����;�W{e%�ß��q�}��ҴgF^ڣ�U���?�\?��j����(밯A�qt�b�Cx��	����R�+g=S�k�S-���m>8H�wr�#=cٕq����Sp�d�3��S]6�d�@;�F��rh���K�9�͊4?��k9�Q��1H]t�k�����c��M��^Ƙ�N�R �U �!j�����'��K�4�}	��a<K����1Yz�&�P)��Se2��]��	�'+z��ꊯ�F�
XZ��܄U����-�q�n�.Y^�4�h���Q�+2��N���	�H�U��얤8p���9_ڎ����b�Mʙq\Q� d�,�N8WW5��o��i�ԀLnճ�u�&�9/�H�|>�#l0K��*��WCP��fR��~�6��.B���N�r"�ED��*>i�-��tC�#���6�FOFo��J?r!�5��Wf����O�È����t(W��Ln��&���f�BM�ͫ����P8�z�K%tS$b�0���;³+`E�Z�]�T��M�/���D�z<��P�3^�)XL��.��+��寪H8]d���%�k��r���[������;�c�66�$�T�l}�@�V�ɀ��P ����V�Ř�Yet}˩�_��]M�s�n�\d	�2������Z j�x�מyy��p��k��J�~�{4n���"Syz+ܸ:|ar}r��j������f��4v�� ���,pQ�G�����C�T#�0r�W�����rÀ6�M����@59�>���$�9I�eےP���b����B��a�K����a��_�$[�����t����T����5����4�*�xb��_���-)?�
hz}��O�d�n=6`·�KE#F�����G佪�/ﶀa`>
WC�~I+JE����u!}:W�!P{Ϣ��D�y��=Y\�Ajj,�f����f ��� �.B�J2�{�96���d�ŵ���ͫ������V�:;��^�N�q��>�w_����i#�L����W��̩_bB�����v�+�0�_���V�踂���u�N���jS��p��c��ϮgǱN�i�b-�҆��D#P,$R���4�9��G�4�S����@�K����0��,v�(��}Iت�70{q��p�k��]�iPq�W��%�� x���y3�~3셑�tq��&��HP�U��l=��P�t�3�q�����X-�p�I_�Y&���'Bc��V�I�ƁUPwfT���i��e]i3w�~� ���h�j�)�<<��
�%9e��aT,^)����A�m4���q"���{�*\�'��wq]���B�7�����.��L/�[�&�Q�4����b�^:�<'��4�v�zcl������dԖ� ��l4\&��s�x#���(���>���J�-jU_(D]����*Kq�)u6e��3�f�$:�s�{��@�$���{�Cʣ����5Z�����a�q�,�ɒuj�}ܨ�����Q�g ta,(�j���e�>
U��O��6���x�����{�j���կ\'�Ka��^��8��-"<� �;��Y0j�H�o.�'O���̕*&�>v�����΅II�����+�p�N^�ِ��u��T������7Nl���9�L�%�`�H��nǊ���e��e�6����a=��F?�tS�;"~��`"M3�[�\}���dpbF�p�פӳ��ե(yn�����Z�B�IgП������ß�r䫭c	�|��9�+�x̓���r�it�P�*��O� m�����-�+��>|�fZ$6�S���[�����_��b���N���~�(_�c[iź�c)�m-�mk��0o��vj*������La�(׆�cX��f��_��E%W�a��P�?�?6�rZ�so��q�HB�t��g#��
c�w.���oԈ�$*�XX���
I��\�)ݕ��g���9y�'���zM�H�Z�Ze~�߂�MI��4f�sct���C�C[8ԅ�dv�d��k�Ƅ&pW�I��!]a��6m�֢�8�|�"YW�" d[ǛARb��N��B~C�qI���@�m�ÍN��:��� z��n]����,F�`�:�=Ԯ֌\��u�f�<���Q�%�h�k}���4�XAA����?�?��@u�@p����=?��΢�>���B.W�6��x;�zn֨�ϗ�u7x�Y�`]9�HEA����G;�0���U�2z���f]�4I���]�~]�^N*_d� umP �M@w�1i�hzNM��ɳ
y#�b'#'/s�D�/4�o�<GK=:pS2?�,�%W:㙲�m�۟g7�}��O��T��t���Ն�;�V��)��9,�kC�������)9���(1���Y�8��T�J�+`�%E/������.��ƪ���m�s����B؝!G�9XtM<�5�6N.?x	A�B}�����Z#�OC9��ΰn�q&T¥��hT�*hX�ǹ�y_�}��U*n��O[���������=�D�z���P�/s�.?fɢث)��i�������ƣ�������+#�7)q8�B{2;�F�~�\���@E1��ǥ�,ro�M�oZ5bJ��U.��T|3��D����b������z^%��Ý��Z�z���oR��f�.a$���>�+@�f��s\�Gx/�Gx�Ns*�N���������_H�1̃���nr�c��Cϓ�V#�0��Z�
���T�X�k�ċ݈3�sY�ٯ��ҽ7/ٗ���p��aޫ��֟u�@\�|��6Q�2���~X -1��SJ�>/�*b���)�t��4�$Z�Z�g.��8K�U�iz?l���T�-�kfi�&;�.�)ݷs���>��:�~D$�+�A�0�񼮼���T
����l��%П��̐Ρ|^n�΢U�DAF�Ŏ��� �H~����������P`2��⑤.�>��1� b�Gn�p��.�kV�q���KD��B8���
��#��s��~����$ntu�Y���c�l����E�*����ov�=�Ϫ�w��n�2��
�/�����D�-;ic��䭱�����<h�4{��\����Ǽ��wUD۰��$Y{p�\�iَ5�/6�ݔ8/�T�S�D�U�"�"i;�Q'F�쩣�'�;��Pv�#͔j.���������DE����ՒK�!��^���a�l�+I�]������c�eo�(t�\ZgU9�XB��*D´Rs��F�-ҽY�����g`��x�.��VOԽ�o�^�MV�)Z)[��Nn���1���rw�����I~F絇��2`��6��:�yuSYu[G�fЛ�	��ڜ�Z1k��R9&jrȺ^�	ۃ�n���A�&'�{�+ψ8<%:��~>(ݗ�_�z��K-���V�PF;��^33�J&��X���2�}�9�ڔ�]���1R!�^��O��#I�zC�RR�ȓ%�ף���X�5�-��1�q3'7r�°p�`����0GL3��[5�P��B�L?st�B�*.X��7q�`��x�1��oG�9���A���P�a�I��V�%7��"4t|6[�c������Уa���H��j��|w��x�Jc>{���$��k���tH)o|j (��v�h6'QW�#���c.Ӹ��Da�F�yr$�k��z84�V��[*l�*��h�נ:�в�.��F�NTHK��x�/w1�Yf�$�!v�H�GC�Z��L��\���M ��ɰ!A2������ZA�5T��Cd�l�{�ֺ������PZc�����ze:�\?�\������%'\-�\ؖή�(i9oVD��r�E�ZR<l�R1CU(��P���Z���:�(�S���-�3�Ϣ���12(,Ң��H�Ji(p����%���^6��
���~�G����Ҁ�^�`D�r�q`�W`��w�se�U�^�5�����Ɂ,5��������<�������5M	x�%j�+��j׾� �;���`�*)�O�d����7|g�Ŋ�f�#	g�~��ri�<R�'B)�\�7��r͆B�wZ�_�Z��0q�u����������NVyBۤd��/�N���g&2K���v/YN�ɪ7��r�ڊ���
��
c��I����i��w�	EN�T �	�B�}�ʭ���^˕)���X�+�4� Y"R{�}r)[@��d��͌��J�;#=�|�F,����ߟh��� �8R!p�
*[���8�����OB���9R1�9����B.��d���.l��v�#	0�k'g`�P��$�`n����{�DI=>0�wGĨF��Cv���2�U>�4�7�y.��z�ý� (���8�4�a��<܇%=�������t������]<�:yV[�4��>7�n�!>���6Q�nLd��%ݎe
AQ r�r�Xߠs��<b.B#���4Ĝ\�n��r��z��ԯA��"�Z��r��e�E��@�ঝ�^��L����6�Z���>:����#��蟌��"MI=���QE��,�F915�r��t	��N@�W����/���(��k��=�<�! y�!�z�p� �&�#��8ђ�Za��P�TZ7r�K0"�"4Ȱ���%P���Z�G1�Z��¦�[X�'��B�N�y0��/9�؍'�:3q)�~�b��MBh-6/�?K�>�lvF��:Lq,0�TENԄT�ZIXGk��d|`�Tph����ЃކQ>�����#)5LZ�|��ɸK1s�'���cC��� &��0�B�#�_Nx���b�(��.WtIF�N�_�k��=e�Has\.���0�J@�w�f�͍��&�'|@�G��snU9��
�nI�_j��!�).VPK��@bz��4sZ��H-�Z;��H6!�wFN�	���Du����N���0.�F�^����ֹ+�����X�B(޳Ç�wv�iWj{���3gi�3S�����:�B�����L�U��$.����C2x��K�ʽO�;p��a�����Eْ��� $ ̐2�#�+
�+s`�,yo�O+���JH}qu��ˤ_�Y��o�ԍI5��|�wl�my��Dȵ P���(Pn�smM��.���Ҳ�G)�*9M��mI�i*?�����i�QKV��
����}��a@�K��#�S�N��/�ܝ���N�C��X{h
�V�<��9b�(.�몾��̵\�3xno7�KC[>*5p�=g��2)�M�H�@��,�������N@���+��'��u�ɏg^�c��*��儞��&�nb�@�iQ�L9�F=?��`�+M����%��d5��<,����ˀ�*l.{�Ou�������*�w;��Ĕ�զ�[��eQݓy�%���g��c~Khl�P�*�b)'���c�v�G�'{�M{�:%��04��ASv����
4$ī��:�c^�`�E��]CuCA~�Ƽ�q��9W��g�xH%���:��Ur�f��Ũ��9�/�^N��Y�5K'���Q7��m����lR��Z�\��vBe~��Q��~�n+G_�&y���X�s��s���>��c��U'�M�a%�?�Io���p�;ɠ�����2���Ѕ(;sH�-#��XL�'8I��B�8�V�_bH�b��J�R>�د~zv�^���4����Ļ2�@K�.��1��t�/���|#-���/�� �xK�F��|,M�+Ů�sK��!�:&�n���`̆yx>��|M%���K;i���W�GW,ٛRY"��`!���B��t�%����>cޘ�KMY�3�ޮ]l�F�	��ҭ"l�9��I}u�'�a/y9랴^������
C�w!����:8y.���5�Ԃ'c5�gt�xG��`�,i��������|d��D¼�^���	�v��b-�P��;���pp��gd�,CI��L}/��\5;������2�E�oVf�<�ض+�Ο�B:���b�i��X��7�-ﲵU�R�1�&,�l];[�Ou��<��e����{�?�Y����&��ꎖ7��C�7tЊ�3���HS��9��WK�OC�:�%w��SqvD�� M3ܚ�#�{�����a��n��^��p�+@C]���H�21�T`�Yk����%Rw�,�7*�`ڌ����� �L��6�e�ȓW�4O%���nB���nR��ɡz�A�dw[��-�m�b�B!�$@oy����0��WL�L���e��ke�q��H�mm��]�(_�,�f��D�<m�`����g�\Uu�l��X���f�����H��
1y�>Z��͙B�,��AǹOsM³���������������|.P\S@
����.6�C��G�	ռ	NC�K�ѽ��6?���V�?�������N�Q�'^cG.�۔L:���H�Nuj�_���9��`��i7�'�B�k���L�_o�)8Gۊ�|9����w��1�>�ƫ��4A��[H+�#�qʻi�a���8��<��E�'2��9D�
Q�Y+��b��Z��ErF�*���#7�Z��<��K�Mn)�g�C�n��
�J��M�ޯ��M�[-�-vɖ�2o���n� �=�-��To$Rt��IƝ��[���j7�!��}�"0����BA��W�{1A����7S�*8�B9�Nf޶��"I��,�+�?��qYH�u��7U��b ��ū�t9*��X{�@�+��FM��΅:���ѺF6p�w�^nX�����g�|<CR��OW�K8��#��_H6;�>l��s����5b����,�@:���jX���w�G��E�&@��I��=1_vOI��x��� v�FܪT�	3��p�:}�
{nj{<�#�^�=Wv�T#�l}rn�+R������ٝf���(
�ܩ�!"��OӔ,������)��Jx�;	�B\6S�ƱH��x�V�ƒ��ѽ,[!.wH����N��2���͞g�Ooݎ_-��6�������3�,8�}�1�c�G�Bq�&��[_U�!�m�Μ�A�� ��q�b���N}a���@+8����Iĺ�pU �
���rE��
xvՎO�V�Q(�����Sl����wr� ѣ�,p���Y�F�ω��2oqʕ������_�'&z����#K�s�i{�~|u�ZB��"���N�x>��~܏uG�].(xש�r��%B�2.��x��~;O�2Jq�*����\�)���R��ޖ%�5[*�H��UN5%�U���\v�`�2^q��@�F�ށ�%P�Ѕ
�L}��;b=���� ����4�pA��%͒�&Ryp�C���K��	��z��+}�|��ra��V8�*�S���)Hy,U�Z�LC~�������s��Gj!/w����*�oT�Q�^sp^��	�&"B��&�:v�tܔ�ʹ�t�2���)�d�BD>x�Ql®�]	����Q �G��~?��v��Q@��{xZ}��W��}�~�t5�i��m�N�~��xr}Ÿ�w������!�z��~Ѕ�t��2���(��{�1@V��J��6��u=���H�p�O��E�8|l����,EK �1�b�]��#�<¶XD4��R�./N�5������>��'���M��ە0�͘��kZH��c�<�&�S����	5)�g	��r�a4ʾ	+�� ��ǎ��X&Bk��J�@߭ѱ9J�\qg���Z���w'i/���a��;�=;/�� Y	��C�
51.�Ky�D�l
��tp�L��$(�~�������M8kةs��)�/�I�����H<5f�+�4�Jd}܍�9�*�/�]�ЉA��%����5{�44]:�~�4ƶk�sS�H���
��^�IuS���&ڑ�3ߣ�7�r����"�� �}*�ޅ��f�w֡@�b��D�3m��BX�N��wJ\a�����LQ����q�-'nA'��?>_+H$g j�V4ܮ6zO������u|!\��K���X�8�XZ�=(W�O"n��U���;��s`����1�瞽�*u!�V�|�ݻ-�9QE	����0�f�?j=����{�ߛ06��3ɵN5/Xo+��ݗe����E��H7� '+��� P���}]p��5gX�, }� �o����^���G������:m	�}� օ)���Ԣ�1Ԋ��a+�Zw���y�W���_�Ų�-L?6ՓX���X��٢��?H�Z�L��-�+���	)+ �
h,&��1Qm�a���9�m�>��x͙8.��n������<fA���8/tx�{�N�㔩9��b���X��qO���-[�I��s=s�ɰ�a�Ll��+��<����#��<>��!�˕C}����~Kp��с��v�Pt�;�����3v�v韦_2�M�����O���͋!���nc�Y(&�E0z��[�܋�kߋYn�B�������:���6b��G�� +����(�8����e���ϊ�Juy����P{��8�>����r��̧������_��a�rn��i g Q���$Xi�+����"�2N�A�B���@�N(�,���LP�.@�|���3�ʥ��Wu���{����=�B��yA�QA����F#�bm4� ���i��mz��o�������<�C�:NW���&O9[Pc�^�z+�d��� u#����p���M���J���	|L~#�Ps��jK�h�N�������,æ�3`�$���wMyI��,(��_4h/�t�����aA"�c�'��&v;�:6�m�] !�ܪ��=g���+	��{CRP���&����w�����A��Ud{cTd[GƟL
�B��� �Œs�ĉV�B?��Qa�*x��{ �b+��YbC.H��X�D��0x;�_ Yp���7��H`8 P�&7�E�:�&r�7]E/�&���ȹ����v�ԿW�:���2�Oɘ��O~����=Ȥ]�E!�F����Ez�����I�G��]�B���E2����j�2��΄�54"0+,���Py?,���RJ�x�ԇ�� Ӫ��3~od�6&�G�\*KJ���vy�R#~�*�%�v�D���#�r>=Ȋ��6��Q��X�7O[H^V����>+Qo��{\���̛� ��oɱR���z�QH����YG���-OT��	��a�ʆx�)H�.y�`^���#`ِm�]���w�l\(͖>Vm[aW ��1KɊ�<���I�|-�
P0�`�
�Fb�R����ߛZ�Ւ�6	�9A��e.�A rt��?C.���fɢ_$�8*G�W���p����
����e�����P��:Va������<O$(]�1��ܺIk���5%�69�̮��9��Oe1;�,����-U��/[��2�Wc�Ŗ��e�"���pq����zb�����wH�=���՜�������M8�@&�����1Ú7�1l���������/j�U�1�;Q�u�]}	���hJ.$���z�qG;!3`�J0����b�j���vOg�f�y�=�`���\�4ƬNi��3�˒紡6k�F#B)N�M������"U��f�K��`@�6}.���CS��T�H��m���q�G� a��1��\�W�:�;ٜ��oስ�����+�}ǩs�̺�$��.z&��a��8HR�A�u7�r���iR�^�5�O��R��r���FTD�@k�7f�z�ػHA����GЄ���M�c½��:T-:'�)H3M2v���]fhkv�r�U0!o����Ts�@?��-�uB!D�w���Do��NF����oE�?�ի�Κ	�X(P����EF~_���LƷ�֏��� #�X5�l�d**T�K4�o�O��F��vI>zh!o.�v�xFw���P�'��F��"1;����XG$�6bK_0S,�0Q�q&m��5΂�ho���Yw�P���*?̧��0�k��P{W��+�����+y@�)��	�x�c&/b�d9X��k�*�]nH�W��˳���D��i���֪��C|):�k�&�{����F���u�[8��_�+#@�
��q�pO�N�Mg �1�y���zZ�<so�)ޙ��������;���~(���2g�H�W`�$pc��&h�^6�\\�Ǖ�ۺyf�ך��nk��"5Т��j�&�f�j׃�~A���w����Ǵ�+���؛3-y7[���r�j���sPp	/�q���X�߶��Oq���g�igŁF��t�~�,�Q�u	�I�?#E�[Bqµ��U�=}�+g#����;�_���Li�#���QŬ��� �Gӵ=
��y1���<Z@\�DjQ��tz>���Ժ�i�+�Ħ�-?p&����a��!��H$i% ��ia�C�j��u>8����ũ(��1N���d��>Q�-Bz���m�	��W�+��%��5'+G�F����g$Էhu��d��]gAT���/�Ҡ�(�K��������jă_�R�>x�n=��A]Q/�fR��N���LR�_%����L����ǃ���o����Pܫ� 6ޖ��۶sl��L
����o"����j��L�|�"%�����X��G���=�R���S4���ҿ[��N�y�璢��޾���y< �ps���r�h�Ju�p=P�q�ך��3��B��'�Yޯ3��������4�c�K5�_
Ҿ�]�O���;�Z�K��ǔ?��Ys�2qD�QHV6ÁfI��Z��Kk��r�W3\֏8�E���/m��j���o�J�&�=�}P^WU$��1h^�裸A3�g����>1Ul��5L����|��b񸻚�p$cD�A�j'��̗'�54�y�u�]�{aq�I��ΰO��odvh "STh]�� ��@�=���Pe
���@��b̠˃�珿��^��v>�͵�R/X��*t4w�F��H"ɉi�]��އ�����H�����)0���F�`�*��ޓ�l$9K� D0"��VҔ��ؓ7�1lOp!��ِ�yF���IN�9H�$=��t���H�`�g��M��*t��|mF\�Ϸ�&��]X!��{Z/��;T��9��v�2q�A������A�d��Tq�X�F�������,�������_��Lk��&�~(��>��/'>B�K��
~X��������2�'�����6�i��jLO<|����j��
*V�G%!$ar<�*���0z����Ьv0�A�u��+�
g��w;ըzX�#��bx{ƒfEy�c�����[s�C�OT7�
�R��Vؤ�!v��MPJǦ���>��x4�?�B��#4����tlc��6�z/A�2� �j���ڱz��"��>��{N�T,MhcH>�m3�|�+%q��Q<�n,H(�9�I��ר9�<pɇH�Q��o��ǿC(q��r�8�;�T������i��,tͰ��i�WV6�B��+n��,s�u���@�q;� �!�r��� ��~��w8X�r � T'�,Ae��I`K�Lf����������"�t�w��傾I�>�R���G���-�Ш��fEf����CZZM��=���4��q.{�%Б�Ɛo�϶��4o�F������A�_Cy��f�-��(d�pz�i��ZF=)�,��R����Mt"� 3�W�T��
��۶u3F�Q]oS�N�s,,M��舖\����I�F���"hT��>FG����@[�Gb�G�G6)/ߍo���z�"Gv'=F���X�0�'U2/�뉪�*E��Յ�t��ە^�U�zy	��7�W�؊b�JLm�3(HE�Kr'���cB�Qt��<H�g��h�7�-n�G�M	`��V	�!%��(��.��Zr7��;@+d�J ���4w���̿�-M����x��OM��ٷ]7�3�����F��挄�yZ��r]��ߵ7-���Snu'$0�3��$n�ũ�u)�q�
�� 
*�]A�*��)����x��$2��d����d��F��V�1L~pdR��`
��n8I � �rk�0�<�
Ő�����]�mh��^5�?E�!��NU�q�ս��H���M���R g5:_�����w�|��*�����C�]:��D���+�=xdo�P�j��$�c��$�rY �2!8�0��y!���E��|	�{����R�s�3ަg_��-\��Z���qm�F�8&ֽ�����,�{�lj=�2�������a���<se�`αbY��i��!^�ϟU�w�U+�_rbE"t;����$O��|8����4چ��x���~,wD�ǑuvT���
���ǄD���9��*6��ʉX+ju��\t0t��]5�J	�
�Q�Scg8�S�3�+��q��Ǖ2�K���C��p���V+tJs�>��Y��&H��u4&��02�i>�%�]�P@��@�;;��ݜ)�U�%+�d��	A7n��䏾w�}QPl������6����םzL���� ��61�K=o���R�O<���:��ڙt�d�B ZLH���C���R f�)�4�����l�>���-CD_��xcò�����9 ��ޱ��y��T[��e�׌�)A,��R�|E#���4���@�Zs]���_�4v���)Ĝ�KeG_S�泀��=m�lH����-�G!L[*�9�^:1\�d΅U���!c�zj��Mܻ��Q�J��� qҔ��ɚb3?�h@C�D�7�qS��{��֣��4;��,x�K�<pϨ{�u���Eh����
�1�
}K�	W{�,���⪀x_�E�OA,��juY�Ǘ�M�>��I�5<��Q�s$`�3���D+��.�+=N0�Rۀ�4,~a�TL4�Y�Gn�o�R���]�i�΂do�_
2?�y�09�D�c&����+#�& Q3��-~��M�*y?u��@u�!��e�mǽ�p�����SB�?��޿�{h�tӧH�ڻ��B<:�ۘ^D�[�y�;ovQ���pā�w�����^����@")�IH�.����RS�D5{�ޔ��;�=�C�}��$CR�-B�J�w.F�����4�>��8ڢd?��I�T�ݱ�=�7"Oߙ��hI�5b�W�w e=dy�7� ��Fa��R�}���w�>!������y��M �̄EO<��������1���BLF1���(1ڔ�����Q�N�4��S�,��0_�k�l}��?�m���F�aEeI7h)6 �d�������9��>3+Z���*���������g7�֬9a������6�]W�%Tx~W�L|p�,�v|�UF�����=���d1��Ye&0?��-��msa�n0W���t�q�y��剺my)U�^0�\Q;��ܯ�=cr������i����l�2�W�|���š<(I�#�ܥ#G��)C�L>pYC;�+>����nļ"�Ɲ.�ҁ�H��|����o]n��U��ix��:� �Ƨ�r�� \?��0ّm�K������������>%���m���t�H�F%�ǘg����4���H�%���;��J�"�|�ʶ�H˫�eH�f�xs��=5��݋�Ow`��i�0���%�{�!��xU�d>��\L��H����<cE�*���gL;B3�Sa�����e4���8�;/����E��5q>?���_bQ�=O��a�q��4$Fa��5���< �O��QG^��_!%P��ɛ�Isz�eaj���cT����Lp���i�g[ku�KY-�6�!V��!��:c�_ʇ���	SS��̤5�m�5�6�����S1��2V����B�L�/�8���Q�R(�ƻ�v+K��Tmݝr?�6��Y5�pAzaŇpH�U��h��(�3��W�\3�ɝ�֯)�܏��P���uu1�=	3���x�!J7