��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%���l��o[��ɴ����>�$��	6������b@�	������b��VJ�o.y����L4���Z��1룠������	�<�~���E`��-�R`��k��-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_d
�t!���N�S��گ/�TNM{�C�5���M��;����L�S�:�{���\p<��)�0W��B�R<Qt��Ԁj,3Ӂ�v��`s�HW��眣�U�Z.͓k����W�z�N��VXi^�p�ޒ�}�7�"�U��J!J2Z�O�.A�u��Ξ���eb,�[��ޞ|���HW���o^�O�Ǆ\:/�"�?c}Z���⺈�7kw;[|X@eA�!*�KU��V�8ߚ�?#�F���񃅭����M3�Og ����O����d�T����qM���\F�B4��Ol���].��W؛r����܋����س������ɬ���3�`�b�=��F�k��jg�\8�D�FON���Q;�(�h����j	�y�����BO�)�܍�V��
d{:~N�fH�O��{��<uD&*���%H�R9�J+o�Q��6�4P�v�8ƞH�o���W#�#��Ϳ���tߠ?*Kz��l'��}ُ�7@@��\�7�K�L]��>6��Ǡ7����� �Mb׏&C�16��Z�l��lc����N�tQ��=��+,�k �:�����6���𝇏�����t׫��Aw�;�V���ly����Mt\���Dk+���l⻬� ��y�Սߪ�����b1},֨|N�Ek���|=��4�"�+���}
pU�R��B��П%4��dG����Vj�l�E���Y�(Gi�Q.�(����=C�]�n�N��_v�k���qmFt�X3Q'Ӽ�j�Zɸ��i�Cw^:�;gՉԯ�M��6�� ��4�
m��%2{�*�Ѡ�Z��j}Q��ܞ������:��>����p)E��/~�8��*9�����T�2�#td��2oÕt�6	�NUu^Y�����;��*����D+ȱ9��IKaU݃�B���L�G�=�d'������� �c�E�5��$%�o[&@�T7����y�z.�u���e��~x���1�D�࿝��~Te��$�Oz+�"��=��O��� ���k���CBL@��ɠ2>�=@��b9ۣ�QҚ�n�E��8I:Nջ:���B���]K��(P��,3ޢ�i}�M��6b6mD�~�H��j��d!o�7���������P0r�+�؅���<M~X$���
g +��A!C��<4�aJC%��f@�B$QRw��:5���~Yਚ�Y�����*��-�N�0��_��t�9.�]���5�����`2�ա���s�N��;Y遼��������g�+}\�)H���jlt�xz1��Z'�9��v!�a�s�9E����[�1[����k�BI�䡝�����\�Cz��4�7JW_:��9(�U��t�����֘��󖭧�N�r!D�����監�l�}�J�?�FY���NtD��C��u+:>�2 ��N9����n�߳���V*�Y�����;�8sy^yv�c#�����s捹/Q#v�e!q�Gz1�Y?~ܛd\��ϻ�T[����]��*�%�~N��QE�"�_5M��{LR>O��z�]o_��Hs"H�(7��&̣��8�C�7�r@6�Ҋ|h�����l��t\.D�rYQC�iB��{P�'�E��F-J���FOM�|�I<��y_��#�:F��?~� ���.��ce�P�!)�����،GR@���2`����g���'�&�Ԗ�c��ǎ���Fﯚ��9�۠�0R���P	���Bba*�h�Ȏ|_��Q<1K�.��-e���k
�(NF0~ך���Q�g[� ��c�{�gq�I�x�$�V�єo��˺(�&�N6�/�e�TO��~���)إW�C��2|V��{f��!*Z�⸌�������8I��z�k)w�}�?}�87�+1�s�����&�8ӆ�J��"u ���H$�?�Z�b	�Z�\*c=����[s�4D���w�Cw�q�v5;oތ��CE~Ϋ�WeO�9{���U��h���v,]�����N����]��V�l���
�h�&Ȣ�ik�̶\8��/�Q�h�و2��M�m`d�7��U��J+淆x�0R\��[�3s#=!�z)q@�A&�O��NiH$���~'�gB���O)�-88�S��w�e/��@�0�ly�_n�F�� ���_�H�GB3LɚQ �"�0����<�W�dTDE�D2B���؋��|����?�e�M$���J���A�ۛؕ�<���ho�P���g�AxL���u��[µޢ�j+(o�O��f�	)1~*~����߄S�i�)M�'�+(��m��\�=],���T\ܖQ[u�"�8j$��#��ԁ}�n�o'v�NxjU���h&���T���yآ�H�ܦ<�Ӄ�;���g_�[W*��>G�� s�#=9�,h�������_���igNg���g�J˸%s&W�v��v�2�Y���lf���bu�����Aj3�9gBY95	�51��_��������;��>m=�eB"(pV�A�`[B��:��7���%7 u4�D�Dyp�`��s�14�$��כ���S�rZ\gr��6΄Y������!��"1�����J��| &DC�ұ~�B�c2{�ܥ裆�(P������u���[4�k�����)=pf�Wi��$���+sl�	P�q�i7�ͶG���L�2�̮�>lnW�Cܧ�S��)���' �ڇ���t��u��'�kQ�Z&�q���x3���)��@��
x��g�[��w��T|����<R�ϓ��F��#�]Z,��!���G�zyǺyћ?�!:>�;�xFIM� �����ö�c�LA��2��&@{LOmI_�ѩ���Y�n"���ܯh���++ַG�8!T��8�m$,[N�ծ�T*;A��A=� ��DN���v��(�e�ຓT9]��(�O���ؙ�#�s����	g���*
-T㊜+��oA�^��`S0#B�5F�7F��c��t��N���2B �'ᶞŵY=uWo6�h.3�u�nj�l,�]dU�����v�(E�;�Jsy�&���X��t�l�U��R�3o���c�;�)@(F�K<6��E�L�����?�N��<[�/��9���~��E���I�3�'�덥�5���S�-���Cc�t��[կX�������p ��'u .kg'�(�����f�;J�4�m
)�W�"n]��ꇊM�(�9Ey_ϥ��e-%o.��A��Km�Qcʉ�%#_��z'7�z�9�g�_��ȎE�u���ֶ�"Qq�Z<��\����ņ��݌���M[��;�є���\�r..8{��}o6?���az:�HrL�ͽN��x��@���N�L�26��9ě�Cz0J@'.�����-Q{S~�Mj!����-���JVه���O�#�b���C�)��ݷ�Y�~��GH1AE_e�È�k�γf��9y`�L�H���y���w��BJ�ħ�%��&�A+�%c�7��-D�TL��ܨw��Ђ/�}�n��4!��̒�:T��z�Ksv�0j�4���^?q���`��@L{�*S��g&^����-}]�����P��7L�,	jQ����3k����;!�+��G\}�îMu`F��,�z�6��FW�L��C�� y'^�np40�">�g�K�9���N�t�;��8�!�-�N�%^e�C����b�IJ�<� �ؓz������8e"8��ĶVP/���uۇ�У�k���>��*�}�{�_�4�M�I'	r[,M��8�z����m�2��Vɥ��9���k�k��O����⫉�M�#��(���ay"��8�A5����($Z�Wxm"u�k¬��pQo��7�r�^ �װZ�ɂ}JF;�Uxi'����Dw1&6OI�Sي��`?�����S�W|�?,R�V�x̨0K@;�
h��*X��A$ei��퐌P�d1�}��z[��Y��ё<�O��K�X-fQ�B�:�5��3��� �n	�K����h�2Q�"u��efx��r�كU@�L0�N�+���(=D��V�"ߴꇑm�t:ҫ),�Z>פA�#WJ'%J�����}5�iv'F��\���w��ôb��	�t�>�U���8�0:��5�g&�D)�����	5=T��.(M�����է��~vRh�syeTz�-	T�0hW:ƞ1�G#ƅc!Cvflf3j�n��������"��o��	;��\��F'�N6�Τ�z�s�N,�x�W��h�^�U�J�����x���Ȏ��:��ӎ�`.w�E�?}�"u��B���B,�UWX"�2�З$'?-3��m%>�M�0�X8�S< V\�_�q 4�m{GTm?����'Y�M���S;�IiBW�|b��t;��&ث���^�:WS��M�P�WF~����	A 5����xHMN,]�z������*H���ٝ!d��$������j�\j;s�~j�B���=�x�""J��Zϋ�Oz"��G��@1q�	Ed�%��6]�6��B^eYꆟ�i�£��x�&! �fC��e�ߔ\��<����I�eLd�d�4R�;ŝ$&<�؍��� F�"kk��
�`�҄(;Z�.AmYDt�.\�Sy�g�
�V���\E.�Y$]�<.��n���暳z�;AB�D~
�P�Z�2�Z}L+�L�45L�d���<�'i��7t���s�nW�-�X[�!�w7
ܴ�^u;+�� �ݪ؈*���Ar㐄R#�O��Ob�	J�[G��j!����F�瞐 �F���	e�������`bԶ���F�®a*���VE�ȩil�����p7��Vt%�k�ɛ�
�"�3�g�֑�0�<9�0X���[�y�wF5��,�������ͨl̢L΁�������1r 5p��WS`�lWژ6�L���5��o�#�[�*w�#b&�a�UwpDM�΁Ø���I��o�a�1.�wBʒ�*X�#�1�v\�R��@�=� x!�x�I���-/�0���,�2��ӵ�I�������o��,�� �W���R��.�ȑ�=V�+B`�ї�	DD.��fq��Q��!]��[�u�?l繩}o�E�s�Y>&`F碁ٵl#��O�)`YnC�E^�XH���%ܤ��)G���M��Q��n�_H��_��ߕ�hl��@xR��~Eǔ���ՙk<! B���~�n�2P'��!�K龃@�*}�:�5�4	1�����`��d��/���K��Q�R�	 ӂ�k�Ӟ��J:��m,W�%�BҀ�y�ZV{�&�>Y�(5�bDţp�THl>�+,�����lo�Ξ_g�K����C��ͤ�c��}���Ϧ!��Q����Ng�g���r����O���cgD:��*f��InǦէ�"��Ь ���W�E	\�emJ�x�e�E�hA��
}�{�H��4���"E'jG���-����rd~��f0 ��$1ץ��E��9���H6�v���dR�^%�(X]�d���+3;A�^��x͛�L7P�L�6|��l���uO��T+e똙��S�f2m�:=�E��(�ǓGp���H���w2NJ�=94�h ���k�i>Xei�S��+�d�����%f�ڏ��N���Έ1��V�s�i��r�z�2-X�E|hbx��դ��54ies����80���7�p|�$�U�~��r�%��-�wDI���;�"���lw�s�����E۝E���Ӏtq�H�dm�r(�]3Q��pG .>�����e;~�*r��d#S�~��Ǜ�_[O�,+!�?N�0�|2��� ����9Čvu���MYA�뎇i�ng���Q��_	�a�'+�!�W��w!4��j�5��A^��QX2��<5�o��C�y&��0�\߷�����ٙ�o��OU���@���r�r���:�i�N����F��Sa;������rl;�j�mG0pq�+p_w��B�R����_[%˥�z��n��J���sL��3/ד����k�꤯��F��J\�l��y�LTޗT�s���}���ep�
e>�������B��h]�u(a�./1��Q�|�����Gp�i�Mf����pM�E�F��y̓����evP\���ʢ��wZ�c� Q��ܺ���pXگ��n����@\�v!��&¢	c�I�ڧ��E�4h�̯�l�mr(�u��v�m[ǠY%�/�Y��+��z������4x��OT���l���-GݦB�̶wV��Bz�T����|�3$�[S�s!�Sī�ﳃ0��ƅ�w��Vg��fRn#v�w�\PF+I7_��w9O- 	uNj�?��v+��N�U�U[m���
묥��X0�6`�e�?�ܲ<c��ZU/�%�\�:H�ԏ/^�,
����Xk1�W9=H�����#�K�}Q�R͖�k��jO+�T��ve3�I,�D�rG�?�cP
2FcG+9:� M�t��A�l?7p���lj������s�NF{&�R��MH�/;�Rj�Q�AI:оE��G�^
�z���~�Z����׿���w�}n�L�4�K����S��M~L,����5�n�%T��7[I���y����|#jiBsW���,odN�=E𩝸|�5���~����k�Ibv��I������fis�g��뚢��{���e�T�ѪT18��b��I'֓��ѽ�>n�v=��F��L�g&iJ���Ӆ����1��4X3akQ9t�!�o[S���:�
�u0:��t8EW9R�t����-"�A�aQ�9�[v�V�
SP�%N����ԯO�˩B���v�ˬ����8QX���G�a�耆��=@쌶{�����[@$�+o�z�y���nS$�sv[���'K/�����"��k�������6�o�4��|M�~��[� S���#�kH*���V�kԽ�׏Ą������j�r��1�t^`���☺�@�Uy�*gc�4�[��ñf�{^kl�ё(KxYD�?��,��}Y�����役
���c6��:Y�R��]��q�B`�?g3D�T�p`���A�u�*�Q�QʠP�C�c{�)I3��sF��5���Y��pf�޻���JlG�&*YG�HL��W\+;K�n��k/\T~���]ٟ��!CN�::�j�,���q�ɏ��5������ŉ�<���u4ݽ=�a�m���p��������f���E	�Wn�>w�q��Ղ���L`e��S�A�p8ڧ�U�s<{���!�ͩ��m�i��J�{ (ڳ���/n��.�f���y�4��[��s���|��`lJ	�`�3�����M�U��o���C��3ȴΙ�s/�9���B����R��b@�n��%��iR�+is��xC�<'A_ms�p�Nv�Ê�]�ޏ�ᨔֵE	��,��Dxrvq~C��S1kVv(��G��� �����j:ي�.^k���g �ֱ-�]Q���<cN�K���q�/��ɘ�	��GJ{M�8�ˉ�*��ImoD>Us;�"���|����BM0���9͓pϏW���_I��u"�hIY���|�Q]U$CX���ne��p���X�����/�3���@)�v��B��p\	థPȣ���N�;> �;��M�Nv��:|��kM�O�����oN���Y���e?�M�,p�Uu�B��c��C�qW��.��4��Y:�T�q5��l����A���c r$Q�Egh>3x����;�!233cxB�`��;G�.#��3Yx�ك�>��R�����׵�%���5�Lr�[���"���4:~5~ӵ&����7n8�:]r0.�K+`��8�:W�u�B�+���w{��'�,���Qa�i�`�Y{���u#�%$0��	�P�RG��C=_� $�)W����wͽ�] 'B^�pg��Z������#�z_>��0�����A>�5EX(�;�?r7�w0Cp�K�< )O��$?=ZҮ�p+z`�r�x��X^`�})<�u�B�1~�Ư�N)�� Қ��Y!�B:��dp�r��p�Ѣc�%a��s��*�(!*M�V�"�0���"�tQ�gڥ�>1"��/�xc��q,PJh�����{��o!�+��-�	����.p)U�mQz8��'a�k�bM�b�������,|f=����}�i�	���^���yl�zk��&zg�h�Bo4�±�Ô�s 1��,�"�j8��+W`-H�D&����$�U���7�@����m��yTM���@���/K�MΚ��m���U�C� �Ί�+�>h�:��!Q}I
Zd�ZWn��s�:	-�;/�!O��ά� AT��/4�	;Ⴒ��N��T�W���z���}��@r����{��A�k��.hMn�V�O�l: ZB:`T�T���^L�j��p>Ъ: ѫ����;�^�,r�rd��u�vmD�c�.�v��Ex���j+�83<�#�����N�	���v�;f�վ��+=B�eS�vU��׸˓��(����򖪦��y�� �E5 8}�*S���*���Ѽ����O����z'e��3{�=#vu7��D�ɿ2Q���k����t%���tL3���n]qޚ\%�R϶�e������H�[�]a�[-��pA ��������a5�����A�,�Q�����KS
��S�'��5(�$#�\���%@�t��{�s�C���3����ۨzz`̏FB4Qr'�)y��M�n4���,�o�b�I`��-�=6�{p���a���y4G���v.�~ݯ�2��|ט]԰��!k�<�%+Ά�&��Ef���������fS'PT�������C��|��%q�|rF��aֺ��K����H��\��xř�C�PFj�i��O�!��<W~G��[t����ڧq���+w�<����?u]U��;��w�ă��i�X��k�wmc��CY�1�;9bZ�u�>�7�{||���s&D0��E��6瘲�@`�=�J_͍�����W�F�2��c�B�n{�^c����؂�R`��+�U���떂a�����[�vڨ�)��bG�=T� ���]�KP)������>\�Fw�b�徾M���h��ݰ��P���7�Z�KM���̚'}�$��?��l�V$����5!�Q��c���z�-J�!.���ص�Nr,��I]����"�H.�)���d&����U!<��F]���S8Y���@�����a�cԆ���.8�xL�$D˓���-�uR�LR�:��t_���=I�t�A��F3���=��������Z@�
��>}H�O`����O�B{̭�t:�؆�7x���ӄZ�mnHvV��nE�~h�D�����me �	���HM�T���F?3������jZCO0�;,�I��j��3ǧ�,�y�ͦ�j�����!��
���o 	7Z��8oxEF}Q�O+�k���#?���ӥ�ͭ�I�_�Ma$����'-4��p�J����S�C�tk8�w�(�O���_f!HK�ܢ���y-/�,�D�*�AT�-A���mKRJ3+�`�'�鄷[���Xɰ��pF	V�k�!m&mL���e�y�AG��0ڗ˘�y���z{��N�H��fU�Zr��I��5H4:�i�q~����'r�(��{�a<��^�G�֞t�j���!勳��iPR�GE4x/RGK����4󚍞�3�6�l�z��R����&�֘�ŤPn	,�����IN@ Π#�>ў�W
��{�ZGv�b�z�ܰTV[�,��]@4��4y��ʾ��w���Va\�!�@�ۊ�K���P��A[� �I���eC��D��>1��T�M;��㼅	��q�aJS�|�h�,w��͡�T���l�r�D��9��.����q'_(Qӕ6�k�o�:��d����>�,$�����X/$L��J����H� �c�7D�O�]�EQ�w�j���!P�lj�h�jCy����I׹?8;��2L.��������Ϥ�B��vRق\B]�=��
}ۂ!�TZX&}R�R�J]+�����c�j�+�1�O������@�����H���g䔕N��]�)K 5c��4�f@�S����)ܦi`|w�P����*�vi=y����V�,��/�[���#�;���0JI�D���X�f�"w��-��R*�BԠ ���	�R<]Ia#�Zh�^&��o*�1{~Ɂj�pP>]���ӵ��d4LC���@z�?p[?��C�2��0��x�ݝ����gd�����#���V*N/�x�����#Yn\�����gNIf�,��S�u�9��:�p <��zx�0�+r̢��GO���W�]'�u|�i���[�-#�+d��l�Bc=(v�#�ҫ6��w�AL<,�D�T����
͌A�����S�����]6C�:z�C�n�������/���.k~;e�3�n��x����B��rN��|!�g1ۼV^ܛm����v�����-�2�fژ���ꥇ[7�'�F4̭�\�[[�ĀW(v�9��$D[��a�D��T#���I�������9$`�<�X���sA�^�+E� M���ד��1�XtKXr�F*4�z���ݜ.>���d,Y�W�Hޟ��'=n ��jSDs^bΧ�r/�޾�."��!*T�ܰ���蔟��0�������1��0��RF�^B`v<-���'�h�B�Ws箮^y�̢Ge�Y�::�Tmu�� T�cu0�B��������V���Rm�f�#�R/���9�A67�VI~���tE��d^@Z{Q�t�W�w���k��2l�C��(�bhIA�q,R`��|ji-x�ϧ����]֢��腧�Hʵ�������+�׃3,,�|Y����.2���;S�����2��<�K� ���VàJz|�u�l�t$U��'v�U�����
;)�:6�&#_�Θ���J���|e1�� :]��U���TΨq�ɚ]���������QkF{j���w G>��Oܽ/P(�q`!i)�\5����X�t�p]�=���̂
��Wi7��y���&�4�%J��V���L�z���89���B %�HȪ�_
2���x�p���g�]+���}R�������s{���"�BWoa�����u&w+�i�ik���Ab�[�8�E����F��6����ii�Hh!�	�a������U�IU��l\��L��n+g��>C}�8(�F������*��Tu�^�C�7��f�	k� ��Y�Z�Sҥߠ�/=Ê$�D�K�S8x�Ձ�p�B,J枕;�����+��O
�ou��5�N����.���CN�7E�@q񿽟d�am1���1�i$e�	zT�Trb?�M�Xry���`<�1�����eh��"ݼ�� ��P�����0�kd�1=I*�'>0�w�,�o.x�S�Z����#������^OT�Lf>�J�ٺD�s2Vxj�����$�B�>Ƽa�Dg�k@�����(�}���������CVi�Rlqy6��&����u�3ml8C}W�Й!J\�њ� ��ݔIh�$�li&R�)��A���郜�̖rݽ6�Y6�����6H�C]�M�S� ��l�f������F����z��fw:�f����@��너���*�����n�9��!ch�~��'��jwѨ�f�vxYr��r�D�7�U�"�9єއ�� �Mh�P�%�E�Z�Ib�	��*�jC�R�����'���`J��/:5�[(��:�`� n�����1�,��=��w�]ۭ~���-A3����S�^�oʐ2 �*��Ǚ-�.c.H��!轂�-V�[>��K��!�7��"��Lt�ơ�����%�<��̅n
S<Q�!/^o_:���p��AKً���I��ġk��lW�燺�I:��OB⬓����ƷU���V5܅wzj�`=HFrAx��H4���
��עn����������0�Rx����
C�w�)�	x�1^��\mFW��e�
��Իo����I��:�鑼�7��z��f��e���4����\��30�\�*�
�RNЈ4�K�[C4�$h�b9a�&OI_��;	.1īWaAy0��9C&�$��C��W6������eFO����5��8t��)���rgh��\ځ�U�m�����E}I+2������ȭq�ϥ�t ��M�3�%��mn�_̾Av�"u�3
٢�� \��Lv�KեkAQ��ԱC/ ��v��{��)�w�d<�(Ԓ��]�Z���E�3RWkn��f�Qϣ�?�%�@u6l�.V���wwY���JQ1cD��k�h�b����Y�1��y�Wn	I�8�,@�d��c�>�N�8��»fbL�:��Ɔ�@d��6E���.�{�v���,�`y?SJ:��ھ��y��"7U����`��=⢼`Z��J� �x��K����}\�RY�#446k�S�>ZGH�T�">��@�G��l��⒯�������C�^Fi&7kd6ѩ�Q����XyѶ��j/I��j�;���^�� <X
 ���[ۙN�6H o��> �KI_�PV��;ܲ�����B�wo(l>�m�&W��0���3M-u�Ԧ�y^K���)"���t����]���pD��i/����7�w7�B]��}����#�å�< L�{�\�_�2���a�#	��+l��wt�їc� ��R=܍A�L_r�6Eks�xI(�n���}),Ƽ��4�&o�(�)�$�Ě#4|\Ub�9
�Ё��LZ�}ݤ�eb������@	/N^Ǉ�͠�.)#x)Q�����=�b@yDR��5�M�ƞ�=�G
՗<rF� .��P�k���b�COQ��T�"=��T��Yc�ŦBW%�t_p_�9�	A�O��9��[�V�*��ty2W�,�b��$�뺿Dl���7-�Jl��e����ɔ���6�WA�d�7X%HY�+N���ŶO�	6Y���!L�6Lu�r,�fZ�pF����NNѶ�"�-Lv^�'�3��]���{�������	�.D�a�IX����5̙,&;z���[�3.GA�Ng�Ux�����606�$��%�6�yB����G��N�2�5?���f@����-�}˿щ���l��1������3y�sd�҉���C�Gp�d�������d����}`L��y~壆�+����Tݶ���W��|Ƥ���w��p�q��LH�n��ҏ�?�?��g�>��\F��b@���f{:(��;g�5���C=$=?��(�uE���w$Wj���w"��L�!l7C��"�_~�Wqހ�Z���$��@O�g��F�J:PM���D�Q���Ց�L��'޶��6�fo���b�-���^�jk�J��	G��S��@��G0e��8�,���������ǎ�5�K~��m�ec�[�Wp�:^v�Zx����9,�������s�b~�c���4��W]ϔo�LuZ$���ZA��2b�j.߷��{y��ޱB�1A�W���ㅥ�H>����yQ�xI��6eMA{���d���
E��{�.�?�������%�ab��l,�vݬ:]C���1b�]�ӯ�A�^"k���E{��Auwr[2� �}Y�b�C$d�sg� ��f1��\�q��.�#��2kZ��|��~b�i�'��P��[Ht�k5�$�]��aν�a�v���iĲ�1T4urpr[����G�@�/������~ڶ�)W_��xˡ)�~�q?S�#�,����i�l�Oٌ~�k(�`*�[��(��/�zd����~��rudDM�W����O��b��Onw����n0!�]�R�;�����D�t�ŕ��
J�9�Y{��͸Ibc�13��Y?�-�����3�3��C�<Z��Q��`�p��Ƿ���9A���j�k�Ɛ����z�(��ʘ��B�3(�=4e�?���Չ�r�
���|P^՘YM+����f�%�i:��1���5j��S@l������V5n���R�����[uv��j��axCkf/d��S\���_���,�+a�Xy�j7ZgvmL������Q�H��9�2��e�U��2��b�\�g�J�����s�I�Z����nV�5���B������Y�)w���w�4���x�l�ݶ�m�{�̧�a�Pa$=`�E_y��G�:Bq�J��g<��5��f����L�lFVRl��K7Ÿ�K`�<��Y6����ѯ؍4;��v�6N��>C����dt��S66A�5��%���-j� ��
N�V�}���8ᳺ=Y��׶r��"�A�P�ߪ*H���D�7"êu��Vފ�'*�G=u��H��طZA��=�8bG��t*�H1tYۛ4��.�����H�m����6��\��]y剛���TQ����$�F
oB'?'���1��YS�43%~WgG5��Q��G��5�,��+:j�rW1��ėǨ��	9m�#�oעk�� M,�\����m;y�+���L�fLߞV���>G;�
�1�byP�����ٰ�s$)0s�W�f0��k
K#}�0����8G�2=��k�w�/��-*M� 5����Z *9��Nơ�it)��P���R�I�}�H'"�I��X�g$	<�3R
l<��uQ�V�(����q%�-*l~�T�[y�X�&�y��P����6�/�}RV��r=�d[�r��<0��@�U�2�)Ig����&�1�[�@�|T��?�1(��d�9O�~�`�k�tP��"=��:�6r�e�����%��p��a�Q�=���z�-(Y��d�襍8�au�P����
Tt���M3��&|�����1p��!�<+��rUD�����1�`�5�S�ٌUnw#�3�%(���!ϩ ֚<R�/��nqd��Q�~bY�	��Ԝc0���&aC��D�w��P�+Zw1ˌ�=�q�%/2�X/�end�L#]��]�ї{��Ÿ|�\?���AI}!��7\�<M��9����!D'u�X�͕�rs'}@��ʧ�����1������������ByKz��n����XYp[$\�����ܬ� i���4%hH\��j�ҩ�����l�V-������XK��"�����Ċ-���V�m�$h�q����cG�+Jf#Ж�h�� [ԧ�ǔ� ��kXfv]@v�?���Zt�Jo�R�����io�������O�@��­��F�5�*Q�ǷtY_}�"8�P(�b�Zd���h#�8�(���,��Y�� �������o�(�k�ghs���L��ۿ_�6����l��Hɽ�W����/���o݅rƘ4�Q�F�'�������jc8��B����p�{ ��*��,o�xu������ֶ�#r������?�������w�֨*��Q��Ӊ?���j�s�F��t��θ7G��M�W8�趝�-�?���%�n�b�"@��T�W��y� �O���o	8�#��n�X3	�E)_3�4g8�[5d�B��M�]tčP�{ ��x�ԉ525���I��.1X[q�a��0��.�#`����S���Տ�<����ݓb�`Pˋ�+Ƿ����v����u�bi�P�GA��o��u5���
�����p9.R0����\Kds�aQ��@�=�%��	x��%���۵_%M�[����@_�;.�k��M��Y��߃�t�ʄ�3L[�� <T�r��>�(I5�y;�)\�Tsu�~!Y<�Kt��1�;�`Ss}牤�
�_��O_����3�''d�>�O?�b���@�0�d�-�*ũ���X�GMCn.xp������F�,{�3K���c�@����~��T�ы���é�_���8^���s�i�L=^��-O�Nf��`N����p���;����mo����?�"�3k+����X��2���L��`�o�����)��͟��rd��Ԥ;��w�MEfr�u2V�>8=��:{��Y��%���A�o,��)��;j,��6|�@�컱1�
�\�ԺcP��Kf;g���d����/�f�$Ɗ �)�8fi/���N?��|��dZ���A�ܰ9��g?lYA�q��N]i�IJ����Jn�ۢ�)��E���kO��Ĺ��٥y��TK/�*��6k�BH.y{nK��>Fr��#F�W���VW �����c���6Ń�G9�En_HB_Ň���:pE�R�'b5&��C�Ka�,��l����%coK�C���[�i�$S`\�k\��1,��-�I�� ��ܚ1;���$����f�}��0�8��lA�\2!ɦ�U#��͠5���	��/����=|c�tD&/o-���퍗{���2�nO}[޸��l��ݠ�,�ѻ4z1��c;h�-��sl��2�A��j���;'>�*��bO���f]rEt��A2à@gs{�"e�&����a���ۄSDS��U������Z�#;T)�h�Y��`����� 2��G@�[g����^��A��@�@����iBmc�37:�]}�V���H|4vWgn�l�=�۸�O�ig^����jE\�#Dj�M��v��85���7ɛ�B��d%��� ���e���u9D��d�s���`��H�,�H��Z�46�
'?[NnQ���U!C�σ���S�����x�J|��E�L �����{�<�q̊͞�U�"�q�4ܙ�R#C�P��z�X3^����X>�%��z��J ఐ�V<�HĎ���˙���3�)�!�l�i����-i�GaY�B�PTz`��6�.U�g�U����7 1���#�'S����a���P~k,����u��UM����;��@d�.E<4�Q���з����=�ƨD��T�i6+��������H5?EM�g4Y�.$�d_�s*A�M����b��Z�t�{ij������!2��=�R �^;��r�R�p��Po�1Bj��	l!D`2
���p��	&���Fޯ���0��W�5���Uc��G��!)p�����x������gZ�	���*��맺�2 ˈ���G7��A$�n̕|�^��V|�;ֶ��2q��t_�d8"��2�ݨ�-�Ɖ�C�DC�����;��OJ�#R����(e� �L-��˘�_��։��െ�#@���O6,0�TH�3�[-�h�v_y�6�(�2jJ��#�шB��y5R����1�?Yi�cuŅ��	+�1k�sC��Y-�x�^a����ߜͪ�iu`+B`e;�[��v)��}�j@��Z����2K_��%T�u�öl��{ۀ��ʵ��C��Y�s]��:Z���p��%4�&��$��ླ�l����i��;$�ߵя�-rh�6�ϖ�g�j����Bn;&�<P��4���0�=L�Ki5�k����՚ �}��t��e�<�����Oc���S���Y�~vP�k���!�!�q��=2T�m3�.i��5t,2h���7:�j"�x^� '�Ԩ�ʌ!:���v#
��޹t/Y�ZK�"|_����4�b1��c��"79�:�AHs�)R��R��G}�������Fh]�I�c'��$m>�6�
�H�e��c��tڷ^��=d4���@��D��V�U4	1-eY4i���L�۰Ez~�z�{E�5޸�aj�)+�bi�h�� �����ײ�QDl�=�ܴ�4�Y]��;��|�P��ϱ���aO��l���zI�n�*a�,(�B��oi��?�n�D �I�D��=X����n��>��If|�*U��Z�@�F*�F�����ʮ5� P����P�ĩ�E�fG��ǎ{�Z@��N�0�C�9�/��@��,{ -�QTŸ�j_�t�e[_�޶LΞp��E
���<�m�,�|:�������r��r������å�אb�lӆ_�µa6>��q@�=��Җ�.�tŅ��o�*�X�/���f���KIڱ�^��Kzp9�m6�|�@���P$>���c,��C�h���H7����IHDA�Ν�����ohwƘХ8�f|p�����|��/�%�=[FmE���}Z�5�
�:�z�vc�]��xd �e�ZLUb�u^�S|�4�^S_ �8#xڏi�$2{���ʶ���m�_�vL�&ҹ����j�O�ZXd��I��):�^@���I~7h�X-}Kb�J�����q�`�
f�����#mq�Z*�~淙ʕ���}#�����|�O��|�d����ӡ�4���v�5���o�c��Տ�w��&[�
�����^�jy����#���)L[�
��Фaa;���xEt�h)1=Ɠ50V�uS؈ѿ��#���*[�^� �ED�L���X(��Ө#�����T�	w�B�y"��,�$d*vO	#�39�ؤ�W���V�
�5..]�? $s����i9�I�;� w���|Z��E���xLj1�g�1$����'�Y�r]�T��r���]}!8��z��X�r�E���Z���;����g4�y���� *P�42o�+��~GI��r�K쨩��7�)^l�u���Z�a�t��J��J2~�I���@��9C�U]��O�%�WC%#չ�C"z�`��Z߱FAx��f��~�����FB�_������~�5���>��=<��Ȇ�cLX0��V;-�vf�����?�$�h�A?� Wm�0�x|;�"�����p�͜ooh���|��PWؽ \^�����Gi/E6�7Ӂ;�̝����l#�C�����Z�-��+$E�jC�������Ӻ�i�;�Wf����b���O4�&ʶY<�fiu ���vJr5�Y�����rd` �����DVE�Z{u��%���d�\��k����e��d�0�����RU"Ybp���o���+�z�T�]��f��U���bq������1�J$����F��q9Y��iWF�
?}V�l��J�g��
���+��AjiF�L8n�*��U�{�8c�����b]O8�		�?ޟj>�RJ���-�b�Rͥ���!�
9�j|����>mmHlJ��>�Z��[82S����Gc!3d7�t�_}��
�B�)�z1�di��x,Zw-�%�n�O�)H[q�1c|7����ɴ����:���x��;�(����
�:*{�!t0|,��1d��<
כ+٬�L&��G�I�G������9�4��������8^����
�s��:9(w������0�/!�T�� ��
��(M��Ue�:	g߹�#�k2H������"���j�O#d�z��0�cm�}�w�Ț�¢�%՗�y�SS��u�?��;�f��"�-�7P�!�m��%
�5�z��Ϊ7�?U���v�Zw��)iY�{Ǯ=m�;�3��\���x��`Q�I-�I����O�w�a������+LҾ�j ]u��Q��������F̂�7���,�)���V������E:"���&��~I�ș[l�/&��:4�\�˓�Q:�\�IkȂ����kƧ���v�1�_o���#Ĕ}e&�7�g,������}���QR�|��t~+z"�j}p��uZշ���Rp�&��b�IzÒ�5�
����SKw��V�1�Q@>�z0T�r�Af;�Ӟ�U�ZR��b. б{"3t����/�� ^��xY�������b�fl�v�'��Y���B��Kԭ��R-�7�r8��8�h���h�	��Q1:�@՛�{N�M�+�K�>c�w[��ф�1��3I*���H�y|���ܩn�y�\��ι�D2d�uߧL��j� Tvb��E�z.�] A"�=��x�.�!7���OX�MDm���M?AS݆Z3ن�c�^�s\�B��� ��u�}$���:O�Rº2p� 4�CN���gw��pP��UUeM�#��6c]�pQ�3`ti�8$D��r�n�Hz�?���N�k�ŻD*���2n�Y�ȏ9��<��$��ÃP�E`��:�H:A��&����g��`�#�!��ΦjS�h2D(�ހ���:�=[�&�/>[W�K���R��{A�iRo����5�"KdsӘ��O;��"�"aw�.����pև\:L�B�H�`E�ND���� �$��>�y欥��R�{����p(�x`���k���5�E�{��L6LM>��=���$�>�#p����{br~�l�^�ؐ�8���SYdR�V��d\����6W���	���`���f��舺�E�Α2��%��}�K��x�BT-9|�����K�D0�?�������	�1�=F\������պ1�����`Qɨ���Wǿ�D�gE=�V���q�?��U������9�+��G�&
�98��
��@�
��)�Oc5L�\��q�!lyO�Bt!y��S��4g�À�9Wi.)%�Q5:��U�'���_��A/K^g�xѶӞ�l�����V�?�͏Dj�Z�m3*k�d!��}}h�����ڡ�6g����%
_�^��!��y�rSӽ*���%���Z4���wiS%��F��8��c�Y�"�K� g:s�"g���'��*�%��~����1_��ܤ������Ǎ�A�X�