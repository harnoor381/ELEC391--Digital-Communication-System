-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
ic2Oyoo1THzXW0/H6orXZBma6GowlB+FUz9hhErK9GkopLCLss8llxgf2GVzvu2IO0c/CPuWNcak
CYn4mx4N8guOXCESy+EMx2HvGgP+fTF/582jZO0KMerJr8IkdRCni/3jBJPl0WI8AioiVlQN9L0Y
u4d52T9o2Cgxtaz1dXH7Jn+NKehG2SyJynmN9AObwgcH0waQ03cifvxWFh42KH6fG3nYoVqBiiFu
cpLug8UvrDcqCGcsb1IkLvQMa7P/fzJiRrSwHqFFc1muUHjbqviCxrfvs32uq23+WFEhWaaP30Pu
vjPwERmeaAc5gmv7qzLT1nUyQCvDCy6pHr+eqw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 39776)
`protect data_block
1Rm8hyyCQR/YOvogeUyPnsj4EaXU6bSdCgmNYlHRKSKxiKgE4ApmE1jv0eweq1hMMv85Pvhc0ij5
f4Uhr1DCYaaCAZsdaujGO4ffVbTmwrmxHKKBWfsxpLgB08sw1uug7s0Crx1pyrPimLhdKoEWD0OE
5oRupqUf5A1FXk2mvU9SFw2Jgr/USoGCsNOw406RmR6NSR/zGdUzvb1t9p9SaQlSA3df1+lJTfB6
8rWpup1Oh1aYN6ISI986q4XpaYHtcuxwhMH+LqgksHUZB9Jbb/jpCsemHRq1dEgHgH43J2843vwT
hTQQG0W9IVlT0CMu5QKmN+ahsesrrfH7LontZm6OnKTrd8QsdhPV/LHACKRkOWmgGDT0haCYnLha
8T5uMRfmDMsn0pBpkt69U1ipbWuNxCPoqIcIv37RO1zZkytMWuy3OtwFhr9plI04caCVVqmdV9Qb
gkSkBispsw5snscyDIGglRyucQJtVi5acZa92yhph3O4JHCdTpMmXLbjDGuytE/hloPYG9sgXUII
hFLed75S+488a/X7jUOw/8KCfeIOJczTCuWkTE7ur0BDSjVlumJ8zfWY57IpJHbZBNY2IhCD4AZ7
MfA4kbv6bBXC/nkpj/Freiej/M17HvzNhqr23ervfa8rHGJDnQq8UJIWSXFMAABmE1u402BJcYkW
Eo8L2F+YeKYp62FMvdWzzhqG0FZ2ekDtuQUpkWr2qkW110qnbHwd4Yq+9jbli/AalGUWCrn3ikOM
bfgKHC7ZZA/8DnKSKxL4Afby6vvgnO2HX5e5MEktbTwExe5mTU+QoAFIJ9YSX02BjxZleRgyfKho
Y0UnTG+hAJcyATyVv36wXbYY1UDubFwO02TfHQ7dIp+noiPRmak5+UYPe7oy4KrWv0/UfmlX7Cq0
UAopE7XlmsPRYngGvfzrwNVR5jedHxTW7OOZun38Ctx+0DlrxMVresDggkbh6COu4hCUmrv9l4XJ
cQs6ZRC4drVC4+DveKNbeJXmtBamJY87R4FcdVFIKC1zYX51bqwtwp9vnS4LcLHgy7j7rQneqjyX
dQexYOb4WazQY3z0EUzul+yu5pF4TwR20iHTl5tMYhiFgjdJlS0t6nY6N5wBszCK0eJlyQkifqNr
qKnFJE0YOiXeMAY73HiUGthIu4VrrHrknwAoYhAKYw2hk6A5CavaxfyDXDekZF3TYJSb3+3IC7US
zkXmkl3QrjbfxZzeRleefafmBN7FgYs3eF9XrHW8hOUWb5MaSDeLGfvCFTKk3nuT8azxxCHJbRQx
FPq7bdvVfDB7SNmQl2PBQzL8K7nH5wz0z2jlxuRVzVOYEfLZ4HtO4Sz8HcUmMrNg+hGqLF2XZB2r
A51RwdPMyyYMnFncLqcOS7f/enw43TqDjyGqk/gaolohKcYz2iA5GHky20GiHaTeS8n429d9QrXT
KqC+M+0MFTaikzuh9UivyvWcbHQ86Iwzu18dQSovHtEQkZwZwBMaVYfsZ3uTUHaQBmHT2DdofwnG
7LDgGHN6ox2lkxQHFNZOu2p8C0A1jjq0/YxoJomjiHMwPqYkk664/IAroMZ9XoAYtOm5l5cOteV/
bKdkuJbTeXlHcINasTGK3BeYCpb39QQqt2qYXP8vvjMgD+QMxBveMZErlhsoMfm8ENtdxRQ3vmgj
63pq+6XK0SApu2p+1lH7WPAiXQ3hzPRth8FDyhsANHGD9rZnNCvSGRpOvWUoFJrusNwMUS4MD96a
LAd7NJcwT81Rb2fJQzCgxyriAOVCYDWIunpPFpIIuNofd4OyryrvBglFiGAJScSBkLVdoN3oGmlg
NxlamcFhMDpQ8ehfJhtTpjoALkFr01azq4N+HvGdDfCHYBv4GIrfIx9SP6MopWpg7vsQnyPBuygg
JSZumDTM+goP8/VEJu7wPJTUFEhMcHHAh2Ljx+f9Q4AH5jBfzcyAgyczWsOfef0Km+cvkTJYce4H
MF1obDAJs4C1rJS3uofHy6gHXxwbtUDsSxWrhDWxSzyn31CVJtq6DAu0oM56ekORL6XFTKN65VP1
0a6mLn5eOgGj6FhlNgSbLVy+2A90AUk+KSkBF2Rt1zLyl2Fmwx0OkJBgirCFxEQQ5Q/KixXI3vsm
yYh0lC9bM+Sv4HzdAce5WSSyDZDLz+9S9rsSWEkSZg+BAOocqA/FB4yAvpAcRwjirF0GxfUZFFY3
7bosDf5teLJfWojBwzvsk3DIkUafQeNfsxtlfs9b5ye1xKRYhnC/F3uqE1rt+KYqaNWt9BRJ8Y02
Ww7oLKQppnEvFcimYwkXDgrw34oMLTsaB4l378H+ujiCPJouXwloS9Tnh7eUxWktVgg8NCNv5MMI
u0rt9mtJLa7sR2A2zQvygEQ9zqaasD8/dPKnEXOPUt+8CBFako08s1EZUZw+GRxFP44GBR+u5XII
8B3fndNwxvjMoTzYRAOF6TjcVts4zDZApEu4VvcAnMPndyxp+PjaE+UvftMw9RyN16zj2eyYMkvk
t5Bb+pO1PcyWq8zGDh0UDHCsvuSK5S/nws2zKPrUSGPBad3xiLZ8TAgy+5bFNpqrAjZ3L7zD2a3j
MNAUmtieIl+4f8f7C40fHTWs8rygSC+QPMPYojRmp02Xg0GW+xwnj0UMwhnkksZtMjX3yxJyElHz
GqJIkRNzRKHLjFZjkQu6hBkJx1a9nWEX9IhsH6rXPNS2Y9AxXscUAH0YKicfjh7vWqKMz7wOwwt6
DO6LoWUvkaam9hAaC67TUqeQxXgbQUDnQ2NkYIymqXPJjdP1PeeWq8ITR4JSLdzYq+2obw/mec9G
nk2Lj1yh7XZS+VDj+9svlY5vS/hp4gnTgIvZlU8LSwYdazYtREwbckqften46qCH58aLAG/wrZME
jdpUk8+piWiMMDFegMYJ74Lj2dTAeiOq42703woDFU8BHNNtYalYdAuE/Loer7bAQlTANDjDwZLT
ebPjlxsBxX6GS5wSUKFfDzpZwolKKWxNFSuJqIQUlLPueHIXS6psH6rC4VrzPU//mPC817ghuqs+
u+szSDpU03q43MbY38qjYG2Kfk8ZIYYXKFwkc/c5aWxQz0MSSiF3U7qJ5RkKiCRYHRRbRDPkTSF8
EEKYBXaD4wCQO16CPYmJU/vbqYhGEKnV9+4xLxuhD24tzUFJloaLL637Jb4ppSBUUoKJYw4IDCt1
cW2kUsLboBNtZ14aiWexh9/3Kf4cUrXY9BGVAVLybVkTlEUDlvOzx0zWt4eThVhDNB/SY36WAQdK
qsTiOdKp39Hf8284fv+66eTGBTSQQAMOgCRtxrj1Np6sOIHaMim7hMFaAxkBacXrcnrJTzY0oltk
cqbHq08y41NGgKvHSDQQZB1GXK+NukvxfOe6XnN0FtDwnbVOPz6eDz6lj15WPT8QoHE+CTdxtSw3
ZMgu6YCL5xfWWiAAoP8nNsFKwd6/tRdf0kjEsDhQpnYSBYRe8wgsNmUScWOI1oLWnunjXlwUNgcd
pVk9MPO6qNJ8tu4PMudUyQA2b/06qvJI3OilWUJSlXL5KP9LhXseI9pnXF+8ck6DJxDBuG28OiOX
OTRCIo3R70ysWivIIcegAfDjNrHlEwPFKDTTH2Bh85hikq9fctHRAH2IcBynIXMKTRFXQivQT0Xs
cXg0jSJWCzxK3v7jDXT7OIIDcSrZ99s52YPh1Btloo3V6WW7HA1u+oMIaAa45MjEwSlpMTOYZ40b
WtFmqNyrlc+oRnrlmsXa66kYmhIicP8F0CcDgPPHvtQ0RVfwKUXhF/K9kocJW6ldFyHfqWuLYkBO
xX+qivQXzjwlEowKed3hLh5SlZEQMNcDzge5jjsNcqD+DGJij/XvIHtx6oWGG+DOm6ELGCsxLbHc
OdTWjZyxjhQvAsSMDBLRRy8p0zMfUb+ooYZzueAdV6XB53TiTLTY9U7WkfNmqkxqxVsdWKh8FDVa
WkOkR8YtSJ9clPK8PA41MxbuHvjbDR7AuGjpK1IkV/hoG8EwnCPunMCiBaKvn4OA9UUc/+pZIgm9
aI8LHPaZnR+Wixyc8hceycsKk+YHdXfnI8w/sg/9QVyWuMpKPceghAptlSkP6cl7dFUG0VFIAajq
hR3kstuPyCUMRaiBL9MVDcAPF3D7ijsj180Oo3//xjMuNkUmywSTufuQxGzTLGynALNZCkU15Bc5
5XSSTZeSxQUflNE1NicbzmhcqWseEN9xd0ZgYRrhTzufQFjXZ2Ud8q1FHwREUenoo6jhneez+/8V
qOpNmrOHvT+ZL6gyMI1noLJWJEKEw3Rke1wEgc2ugfCs8dxESbKki8GWpjwMxWADZAWxzfXqBlm9
m4FtR+LDuWyvwLeGVajgaVPY3VvKq0+8lBBYQZ1qhvHkjCQmmjX8pCdGFIHBDIwvl7LZet4625z8
ELxqhCHnB6FXAH44b/fDzv0KB9G0KZVC9gOP+wpJ/9Xyy5xgXHtmNH25MaAJGfZDLWf09hnKITlr
zYwqfhy3gPcj0/+1pG2U14OwbChbd6zeHFlJAzO2iHUoXgZ9fVLyMNqRTch/XBSYTm0EJRZGSXrg
QIUkcEDKYRiJeMUnjSePZGldmwgzMAVvpDc/SONT3AHRDJD5ZCaLll7aipFOunvvolqgkuMLT6+k
M4GdFtXpy+phoPA1hu32bX4XTdWmLE4S8nSH0NPtyvxBcWbdVlWR48ZZ9Zrauj1fUg6yPY/p559t
Pyu912uiVaS9Z0sT/XSV3taLONmDxYqvxi4wojSJmcyz5Id4pYV8f1Z/2uDfMOUeDd2MU/9QWmxn
1i7S3ZkxB9sBs/JTQKtSXanoezAHI6oh19FEgKvoM6HIa955QmZULrQLp2akvHXusxbNTxQtYNFO
kPAulSia99wFVuq/3fJoc0ufS0wPuwEx5AdFhthHu1ogZ7DSTS/JzNKwAd47HiIpAPyqlYPv5V3X
TEb2QgwQ+UAA15V1rYS1FEPXGPUB2lN+lVr/X6vZpmXcDSnB0yNU5oj0RemaPk9NN7JKmFnnUdjC
iEjrVqVq5scw0I0Gkk80P33e97iHPYJzMv1GrWPY29zF0iIXBGqn2oHv0z1bkLRHl7HMMArSeKhf
ww2NlHI0CnZFA8zJJVD4LomIgjh1tnV5euAUoWqpQxSWZTcLRiR71mDeMvwj547f8j1mCM8CzBHR
6eOXl9IQMcRUu4jl4VhhIimxhvC0mVUPZ00mGbSJys/Zgpe6eiP98Z1MEmQ6QAG60Mimu4dCkX+/
Ph9Zk4g7G6nYxZmBoaH3cCSeOJLz2UEPEufUoLdVQ/hmz22PZikuxZAi7rXzCnQp/y6bZrBZgMUe
fAQ0p6rgpbW5u/QmfF11Ba59yNNmWSUJ38obzjyje9y+09e5rwgRfe9WzEMqNQCErdnylzN0GU1Q
ZWwq6NHlOJbDi7HXukOZYUmJpCf6PPOfS4GG3aq3w9MX4NR4bDCFvMJ7uUYufp9xWgjiCkX2qgFt
vfX0OaTUQ/QqbJj6AEjWIcqyh8ZFWg0wie9vAnoe5krdY6v0F7B1aAj0mfkGEBgbHYrhULNIEajo
0o1otsnlBG6S1nl5TySOA5hNenal7vunaW8YWP+rAHWPXruWGFvV3AoTNjeNckAn9BiYrd1xFDQ8
RJmX300zvkKLRfM/+VUIwhpWbtHvee7db6eMZhZut2HhX9PFtrjd3x4rLYhaldZZ5xDzPHVA4wq/
Z3fCEsWQ/lBti33Mk2akfsNmxuAdGOIGT6F5Ricxbb9kRxRhAaaOEDWPh/wXTH002+A9V2axgfTJ
kXgwNYcCd9+ZeXtpMgEzhp98bJAidH3LuVLz1NCNPMCfbfQZGd7DJgn0VJ9N7HUtKUFyl7lDHjSy
jOP/kPvA6cEufQROjDLjEdSyQzoQCOwYvxCCcK4d/bvuru2sPK677TnoH+cU3P3BdKRN2Hh54REs
8xABbQV9tci7XkFyZCOKXb/kRONI8J8qBZLONFg6RZFVgPJKSQB0zwwU736w01yifEy2fyjAbLb7
6wYeGv4W2miCnLYLiEe7PiEIfK0BuWwy7E7s4Y4FTuHxTi2F87Sp2oHGj9bbcJadLH5Vsn9wqoPM
ArB+EZ269PWc8fxC7koAibR5XAxNoR4BF0mhQZa5BG2f0mJlDStKGdC8/T8Cu4qYZhDFLmt9zpPy
AU4ZRU2GaSlmuLfjZC7u9c3YixKVU5e8Y0BVuEhGEohIOjuR/HdkLEWvU+yIHf0Ex6qZ/6J7uJ9Q
Lm2b0pdCdBam7n7VdP2Kkjgj3xc/wamH2Cq6AD3VX2B2jbtL0V7Iv64siwphi/lzQCK401R5rwMS
RgDjHJepqkjMPfyKgjH/gMJMuvJH7jnxWD/umBwZnCWwS6h00k4h/XsSFm+lsMG11zDhul9PmNcg
1YcipEuzIDfWKKHU/xtGPCYsWtWrSmMjoUlfgc+fhqQCJN6PtEAuP8jq9PYL1KbSAgaRoRPfEJ6O
SrLsaDSRKdcSrWTkSi++rgAo+HrLzkzMx/QlxTQXT9iz7AsJf7Uv6dcJaTEt+JylfodEIA41yRqd
qhevmFFzfv2aq3l2D08uTVWk5CEgze6ePBpacbrX3NxvkvEntei9pIIvjsec7EtNvO3YEYF0ke1I
6HVjBwqzPzBFBZ3zYS9lAc3TsYgrUPb5OljY0GlpvGL8U4kbpvNiQl3onjTG/bNFBJLKlyDuMEOT
y5kf2In2/UHTUTxmNldTOt3TlgTCxXjRS/6q5v0ZC/X3NbAC5AFoLjPipFUO7NWTnlnzyZAoGDWq
N0aAj+pxDmUP92SnH7VCYGHttwlRS6hDBLLVb3TFhiZMIdXojTSEETdNdezjsEYqQHYhD77ffJ7n
Yf2D5niP4mcUzst5uKAkBP9DktOkyOwqRtufqRT/WMyFhedBkYihrucMRmBJJ3kyeTt9+aZ+R9Q5
0BwgUbspqJtxjSnrjoJ8jX2AXaFke1BLniaxkGNXNfUwIAVz87jdV0El6tgsPe9xQ3PC4uM0anml
N8A071EthTBi9OecalO19Z3j6VZMsrH+WZrzRKnT8tkP0f/RFoPw5q+WkrfZv0/hu4hO+C4MSsS7
lnkl82NnwbPl6fw5RcAc2WoUwKcyiClrV+OeFAvpGtvhy71SEbUiVh1OwRTF1Vxwp/pPsLvA/B+A
q9If/p6L1Ww+mkuR1TpxRaiRDgoADRznO+8/sHl5ncLLDw72vksWQ4Y1o1tnl4SNhYPPEy2xVCm6
iwjtlUXfMOAzG9oxrqf5Dbx2TkvXqKpKz2Bxy/5OGGKy37r8zvXo/L3tAs+XZF8Qf+YVDtoYrezI
br4HKwP4xi/9GVUD6Kl59MvhYqopm3Z7Tbxa18qr/BTwhtNODsvI1tKYk2QuYzO74U2SsEY8rR7O
7AAWURn8oBU/cQgNvgxE4Jw7uJ1BgIBrQ4tX7p6oHnFbZhOhURXtAPsbXVpFx7KVD95/y8T3IpXF
Z25dNzFHBc2XyMobpqRMlzIcg2xlJxq4xEWQ8PvMin38E1ZJWKjDDhssJVNIzb3rGUkGgc/wm0zx
nhxpwex7s38ksCe1hgapE2FBRB47FPhMm2lxEcODrz14Y5VjWI9MtBNQipPe9chzURv0I4Cw3H56
beOpQ2W+rbrniJYTtQYFY4DlFidxNK2x3sDjxYjceByc85LaePOBpZ1r2NpKdFTwunTX1lDnEVvW
JIDdZ8Ds+55xgsno7e6Ae/momj/rK/biGG9o5iOHlWX6Gakp1A2pheTpWfXdHNed+/i6FVdU11eq
F091VTu28rK8pM/K6kGR0kz/8SOOkPG1LYI0rhsdbc9t8OnM0ICsTFPa7TLqAULFh5v+0v+SE8+E
Byx+pO0QW1h29G/voGvdRC3AJG0tRFN1kUSZp5NS9fAzdjnexn8LVKoiTJklbQNt4ar+gBK9Hqk7
k64MBewkwxS8HLWdlvg9k3MBASwoSFulZ76MMB+1gJT68mwYuegIS//a+JOMC6vvMK5wCOuMHK3K
gfew60n+929n2ZuuPRU4EObz0byl4s2Q2BURVP3LH8S08X3d4GDx3HE+6nZ4DuwlWx8hhfr0xw0c
3zvXiQTeGa2VObLRf5bLUdeaf1LQHVhyqA7Tw86c6l7z9bB+/jmwZt3G2Ak1bIQVSKwfCTXYGqVO
jX9bHQB/1faPhNf/pWEGQVCO4F5pgMxhsf5AupO7V47JzKfbLeNQ+O5hwQz5arEfJpqZyq84AJB8
Muk1x/KGCZsxffOYUGAZRxfPSgzmAJeAczBAr9xlbXUzyJjjPFg7OfB/tFWEsqpCC+PPjmwYtf5H
AIlVK+pDW2zSVzKsvAGIlsj3oGwO5/XRBvkWAUYGpwoANyjUgaSMk0Q1M591iEIUKFzxHgaDM5Zt
Geowtfst0frV7saTs4PligRMi6uQkw8nqVg8S8vc2IiuLYjKLbcAuv21BqRfvUNDqtXjIeJ6g8PQ
buA3/IKlKRoE+PV+UhzmZwx+hyOVYuwC2McwM4N4gaFuOPKJ6GBqgtv5Xnf26lWKJCV7TajEu69D
s2Tso2D+P1p2L5PTQ5BOSshk5wNLOoUv22oDAVMiLqBQVmnAj3hnrZSenLesvN4Dd5uNUzjEMQIY
lAjqrpzZdrt3GkWeJ8ebJ7IT7v+mzMMEs3Yj19LrUtJL/pW0vqG/M1ePGBG+0U8/Fk+NLv3JgqLL
aleKoa+3rjpKEd2ODLNI5JZdz49lGY2+cMV/sVAVoq1rhIEhObXVts3d3ernNcfnyXKaQz90hWEI
TE/6aH1tBDC5qt1ONBm8CA8n5YkDMtyBKSEi3NAtm9dHxTfSZdrQISWdd9hmZuaXa7LMqQbt74uo
bHuX0U+jLFfCYFlDKJbNm56pgX8iG4vxt3EmIosUxbmq5gYElLkHRNfHxjde+tz8iY4kVo8bvqAE
harXbubhcHA7BLqmH8MArlw9w225rr9tbQePfPtwPb5syricMh73rU2OU+SYU5WyzCb5Fjn+qLm6
gRb5KNQ9vtDjqPQg4XUZmkCzMzmt8KfJX+2VusYrwWQDqRqfEFvFAesxYjnemK3j+Q+ZsD4kARuN
7p5RoxKHzU3K+ttkWMw7C3oj6ocB2ZZwz7Q4xqWhBcxDnoH2HK6ZI2U/l0WPryjKqJN6B3MGiAY3
NFzcBuxoFV8J29NBc1/AvrhuUT/ACrGeJmGUtGjJwgJ2QYwpopeUW4tjvBFUysDkXaLThMGi2OST
qSCnSp5AThZ8zfQUnzB9FCrGb439fnrLvVXE7+Wpx88IB/koczmozw83IR+XLEMlygA8aXxvQMk6
tIpvUMsudhakhhOgYMD38KQPMzmkQb/nkJhrEmHh1sSi1ODlBvtVYnT3MXWdaaq94KrOsLrbuUAc
GTD09t3pOJ3DCerGzHf1xBIVpIASGYvyatgF4bcRtb5rHKy4RUN2veYP+66JUibyWwrs3YQrnndc
uZkNFVY9wyQy2otabACOlshXuLiPQnwJlZacL1jXITzYMBnLhXXE5PfaVhu+2di2HDhUc7JYacNz
qM/xVD2p+Vt0Q6XiwFoUF8G4lnOzQDEP7SRyc3rC/WFGeZDZDS2sUjjh+HnJXO+3QpwSirU571B4
WqKTNy67c/yHqPnu4S/Ui2MuBjOzfc+b9pxA2pLAyGeEXVgOoz+nMh/8C3a3ohWPVUipkKJb4SJo
c1gyxUdlMdwe7Mo+LVhf+NkWBS2zD+h8V85qmuTq+A77seoi8/qFHFG5iGsIf8OVqrgi+H5jLz/x
pEtGa9iusasVyFwcO8b7nptysltnSsLhgBrpMGv7YUK54CgPiU559yo2hlSsw0m6j4JYvZTV7B2p
/BFPZFaSAjP1W+aq4QzSj32DS8T0n513OjfB9StFN/bP9MOYLXYDockRT8j6oVGsJL6XMtBHsHUe
He0Hnva3elkpOZh8q+2QMIo9dTQT/3V47KpkayR74pChjchmepwpqnVc5/N1K1zrOL67xHtw6yOg
scyYbi70cGp687INNtIfZCBEv38+8YTuKSRK3wUF84TESs4hX7sFBbD+k3rg6YEtJt5h9DxqvaE5
I0vNDpZj7ImERhc9thQJKRJsGvPz8xewCTS1bHLgLQefz2+8Pd7t6c0pmTJJmp/jGdJ3JM1AJ8uM
hel8MJNn8oFukSMAEyJr5jGWM4BnusNz2mMA4dLnyPKx7tWGAcjoxyLiTeYet/VvXuBwuj/TO5CQ
rgk+AkVB7xcmWsggrZ+vHBmujWH8HHvGW745NPC5dq39va/PL8fYF8tJ/BcwdcCycBJOOTDTCLXM
oCVxrOY08mvJtazinS3SAKkd20bfOUbzIMxm6woVgzvICbQFkIyvLZhCtOoPUDDyq24E+wmRaig6
w1xqP9PW/TgEh1J38qPoPp9gN34KbAJhJWjuhGVErsVfOrYdo1r24aX48KUnnHh31DnH/dXZRyPD
2aUDGIkZAsOuMTcsh84/kD3cRuMvO7L94GKIi0BO97GdbSbu87LHczPtQJG9LGulxPpPtGJiL52N
81z4Aj6BW+oUlEdgec8zFqbRFLhinOPQh0HBvstqdIF7Ab292nxrOKKMH8MM5SijQRfXjwTHZol+
d3oMX7ON7+MrDTrFaAhaYbEj6E3Z9AsdReeY5AvrK1BUGE4QEWXRIVVcQvY1NstMFW8d3l2hVTCm
vKOlllztIKRdbAYUQhMYrMOyOjQvQHjWpKa48XPOp3Rzt9uycS8/NI5NVwUWc1bqSClSvyztJOOV
bJkLdXN702nyHtB+kwLz00oUe5FEli3Ud3GB9RX/lTXUZx+/UN58Az4bTfIOgls4r3vzi3nCjigm
5EpPeUTm/uWCZOkmGQkNWzXUSk++SadGnWX6INYK19U8ErRadEN6a2jKhRawVsuGTxUqlLG0lzLv
VxIzHRQ8J/JoiGX1jnlQGiuSYuUR27ukebTVhuGWhAYg8dybjlA0ngxe5Lps4N68eoR1+MUBjue+
Pl19gFsGfZpAsSNTL3nJVKQO097dwALAYmWVZWZCRc94+AGTnwiKGj2ZZkNmK870MnVNe2HMkvJl
w1/6LbInNemqfYOV9tY+LkoMj5NnrkkzUNBqtA5Puk0hyFJM9puSHaWz+Z40wU/F/wZ8rT/qnSCd
yPBtDgnCsuXWJJ28BVaX84Ecs/Q9pADKYxZK7SceQqw569uRIch9zXuNHKOkw7yr9kzFSHIo+RkF
zkma3zkhK8ba+pNMBkLbkm6WL/AdvE/jHfbktj+wCkp8LA5iARHMde9pZQ6zQgRNMy18jVJHrFb6
zTpsA2RMObnqiArmmSYSz/yHgdP4EuTXNUnQ2RgH5f0Pye0uDysri72mQbi/o+mQBSX9CPT4hT9i
RVRa5FpSa/YHBuPMNb2P2K4Fii87b9zERCxssepbT3e2QpMZtlmb9T59oETRwEDiQQGRdWJaLlux
ATuE2sB18p7pDT7JF+SSYrfGOc+KOT0mC4gzLqP9+19fTEt+04yns9n0C6mgphVtHDeHYXMS7f9o
EYKQB/TxfnbOV8RBtehfyv8ZXL7d95GHjCliTeMbKgKcCRiin8U8L5ltaboWNr1xeX9A+t8VARxz
r9bHRhCPgmxUIn0PcpasTnADrEG6tZSNKEYdeb6vmPAGkcRCJE7puKcAo7i6Ef0L2Hq8WEhmAWZn
ExY1douGjCt9FPV/ykGq06siiZGWIFOUzim9SHKL8XrE/jyGNbQB/z1O2j3lzzss74/p4AY6cVdD
51H6GWViIxQQu2oGk2PwQVZdM2tPB9l1OXOXmVsqHI9CbkbvZPQiKczjoD1hNeJMbOfX5pM+Ukj8
Lc47lHPAGUwx51pWNetnm5u6JQrq3lZqezzfuzg9beMCrgY7rMuTMWisQ6EA4IPrqPIHb/4rTWGN
av8L/LwX6+j9o3bzQtV6qkY/z4w0wJTl9g0LBkEKVlZGNkytJbF4Bdl79mzpRg3wmMddWLLCyhUz
Kv78SJF96BBTsjKKz+d9Ku6fiF/BwRJ0gCXDq6yxD6V7yotbN8RD/MHrKy+Qfi6F02ZL1A75vq6h
wMf2NWUJtLDoMEGNuDozlEI9GbNSTt2Bl/t6hb/LwGec3d6okL453CC1/4eJpMQB71PSfSZjP1Ea
Am6iPYE7R7n8ORWuCkxhDuWKT9eeQnQw+uh6cpOwQ4XI5YZ0d2qyrewwus4peUAD3sgy+JG7vpMk
Qw393KCh6PftrQz0cKqdVF54C7sYY0L5PVklgLSxUucTB3XW28fEmoOtocS/rgjIC/EquZfhC9KG
DM96pqU/p5C5Jq4wT7RMrzMIVzzoFPDKM5IvHTXN9bd7V+/MA74EqiFskHF5q2Rr/wKcH8lFDZOw
Ui1zndIvHU2VAJN1dg3xUDgxJbNFR4C97Q1fNlanyX3CkFVltZ9mvoJNZDUoPh2/LNRgee0FYrj1
YdMLlFOKCSdH7gYbfAVNwF5qj2vy/ZSISyJN6MyoUKfyh6+KIfCAEHwpxLX1iLUB+GrE1PyPBPyO
wELPhL/nFHdzXQGMEAhA/RmEVo50gX8kNBuNJnWFysmWhLpYXDWzowgpb02wDOO74JspIqJrrz+g
jFyykowMPPFOEpjRBC/d1A6N/czgfwrjLKzkChqult/8DcgemK8f3ReCPDjopEJzTAzqBhN9htW+
dKr82La+Fxsne6qZxZz2ej5LxwSlx/pquDFTFD/S24UuYvAGOT/kIciJVdDCEpHrU5t5YO+iDM4w
Pqsp26+vYEQTnI1mC2S2Xl8rIKUJw6kOIVWiXy5FymAuXEMN00ZL9OUyYnmQ5LLaVt5tAdN4sFvr
gj5VQ6dSi+vlQIpjlbASiG+PfkfF567atbM59UgvITf3a/F50szArDH9+s/fg1/nn5mx2cIMqFOu
5r6bFsv0axzmMFZyJ/OtthTps4QpNsOO67bOPVmlUSQ+nCN0GfstvmXBJmkdl/yCN7V/9kOuL5Fg
ZpI1Er2CTKcI68wMZ5+cFYliarjcbTU/S7Rul2q6n6IOk3rGf/fZFqjXxjWcHRw7Vet0++9KP5zW
ttAqWVtKq0XWEPlVgBexCK6NvBnKwm36E5Wtt2RkCABBIosHq3prtWDHMwPiV7INOYM6129D5rbd
dtPjq1tBn4CntyauuVuV+kfE7YwsxjzmGAeFOykDaZedksBOmWUI2JANaVtuMnSk5gSpBdlMCppg
/FLT4CNf0U495PTxoGnn/bQZ/WOScoC1VSJMvbyE/eL5pUHzjXa3S4sO4lg1zEEGOnUSMpQIQSjU
RPYdby+LKjJSDdEfvngMzdCoyig2ZUU3JUj7cQCK7e7MoxRto00CwoyNolRNoGTYALpSJ4StAM0G
fCDF3zefhogBGC9dLQaYBHfiHTliFS5IDC41iE7TAJ3l3olz11pv0oDLb02CfpU+wWmGS8A6MNht
UujQ5iTRtMT8he8YqvcVW/gbeI1UougnVNaTYQiBcQePsAHrOevFkP90us9goSTnLlQKZzlEFwpD
tN81mgd9tiYS3JG9iI5Key5v4cWB85gScF979r+5xQNn1B8T5w6ZOmBJQPShFkqbl9YMBl9Be7zL
A2Esy0k8aGEAc1GqrJs6+PQp81GfBxu3iCVppS7b7p/tk7OpJxOtfcjlHQhb+V2cWR9Jj2rAFZNb
R9Lcy0y41a4yHIOG/UC+6qXNT/JmSqVrDWXFQJmBJObw6PNkmh07ZzwXD2Pm6Nw0OOuhmr0h3DdL
8SorWLzREEvP11K7XM9sLfxcIVr8kAZqufYnVjGpwMZtIx/I5pv8VnIjMSVv3N8mqrraJHDdTuJp
MhPegiGkd9wUOemfVvyuK66B4OJ9mJ8TRQMtyVQfkjTXdqSxirc8xpeRS/xpTquUW2JV+EvcD7t5
svh0SXxBIBvz4WNujhMJk0kCNc5hJ4TVE+K2kxBlQmxWp8zv3QD9JEXszSwFXjKU7Xet879qRXWz
xWM3OP+fyw4XsTrIZxLArih9QSdDBxZ2CgJReWz9rpC98QOrTKQXZo/kluif0Ibt76L+aRUhogeH
qSKHVdxLTdxwcK9D0dN+PNUL1BNVDzc1npkGTEFpRS6jglR7/m4yvjD7/6nSCPy1UyqXneRK4kT3
xKrCp6wtBO4YzQ/UTVKOZHSqgLDImPXRe2s2mVjrkLzjYud8sY4vnYFyiKfUdoT1RR1Xpsq90uV7
X32074TqA2JXZv0LNf7xQm1mCv4uRSt9sk3OGdYNkIXZ7MWRyTGTjYbLt8ystOegbNwOikKmNrGt
eu2QUhM0o6IYQxcxMvkjTt+eXQUZqEIWGUuzyvgkwkctIEO/SRMiZ1O055HUZBMfzc2GQxp/s46o
RKC8TmJK01CQWZkr6OIRFTuBLPD4LRgkhsdIfQ0wWuV7t7/dGAuEX8rC9JFORQT9QqdNQ6B9k9T2
kTiBe8q0KpTOeLegEJiSs81k91FeZKfMf5I09cKC9OpsqiTdqmyq+xAGlN7JR3zbdMwmhaLIU4Mu
LM5l/b3QmDyDjBo/ZLB8Ntn1SHl0YuBWj+M5udm/wtjyhPB/5MdZQTRql6KsSaQibK3bSSKAUQcV
jJmlxWAbcJ5R3XsAHQOPEb9kawUyWiGk8psYU82llrwlB4IoPtyyr2OCvIVQF/UOQ7p+gK+8F/bj
csnK585vF4gdsOX5/rWxp2s0ZD7blTwEl2AJJt22L5K4wVChDGpB5w3nOWo/00mtaNQLSQA0v9a0
EXeUUmRP0+r0y5vpv3DhEH9QZEPsSy7x4j2dujIdOI1D+V//y4WHITedRBK9Fsr74KERs0c7zhEM
LpqpFVPuWPztaRqee+LECmwc7T422xyZrhb+wi4s/G5zCpXOTd3DRX2r7yhNMyViSqlB6p7192d9
M/7r+WfRcVxo0iVs+mLnq/a+62/i6UmiSKIOulLPVXtNY7r92KhHoYZ5GQc3b1aaMNStdGrkdmAh
s2y1f8ubv8xZIJIcfxm3ekLk8PliK4g9qvxm6XvKRFsLt0JvJmve1om5a+oFUDAHi3TOCe4pWf3m
z7KBjREk7OHfsfPOvmDa2TR+AlPozpi5xmsQ4sZlnYlMrS2tU07MSzyWmaqzPMzjYrUcId8Or1uv
vD/rmYBWkk7d47C03Y5FhyzqphKLmDaAZyKjzEE74csFYSpAKBpqZpbDx09F4S/LTeMdObgEXuwg
Z+0Gxw1qSo8nNShHs/S+eZOnwmoBF3Ml4CKQMuuwRQVnPGL5ldovxvJl2QtxD3qO8e4YVntwvnpy
3yjhGN6sBcELCpOWvDhTshgpQez1VmrUNzLtDMvrhsrHS7Gr6dUshvLtRA+SOx61Vj5OEUXIASs0
wPmpecuYX+JWvk/v+wE5Nk1Y7v3jMnSL70j6Dw12LimYEWzWfx2Ym5ZOgmFercBAZD1a+bPBBf2/
Y6qw1Fn07OL6ANrGrgvCLI0ZZ7sawjERsvavzKpV8UButhfOkR4Nyp9cxr87JBUAYN+4ME30u9Hk
0K+u2EDfKBZzSCpamk9k/E2rlV2ffaKN/fwXNK/wH3nyug7g6etRhdKKy7mjpxunhuz3r2MjEfwg
/Flwa4dXyn5rwIi5HT68/TjG2lSt8DEFOADbC8CWLM80nZZvp4n+CcjLcpMjwxXwQAzpIU4mAMI2
onNG3tC32VksUPKqSKm6uMeMDAs3jY1XadI6dpBV7IxKI7W6PUa/JAQ+pHSlan8D6Hel81RZubxF
IY8Tf+beBWrwECuvC12E/RT4glkjCb1CmY3B5c0xczHSecrR2NUv+YspGuv6ii3mhFG9M/VBPAf7
pqrxUrVrEOn3aHru2DVTTjA3LCfO6Txwt9gsZAD7msNy1ZTqS2rlCEYWVEl5JZa8BvodMn7JllcU
8wEmr8AKhbZGWn2APXUQoDwKoJ6u3xkrb/K3RQRn+yY2WtzysO1P7EFluYlfyO3V132aUwRii1LO
rom5Q0KVvRLwEEltXj9UmNdi9oqr2MwNHL57IowzaiJLLUTFmEfJc5Dd0+CQz0SZNWVYuP/nudIT
O5sPFM0XLsOgMe2H6oSnFmGKIGTXYxwhtN2wMBr7yClK1QFse4DHecf+2U0PncDOiZ8yIVKSunCx
jMGHUKUIK3vg80FHqnj407BQVzPYeCqhD+wAj05rQjmll8LEJV1MJKzqf/jqdu54OBmZMvPhqm1b
s/Ractbis5AuQa/RtjmakAS77QCjLdRd9nAfPHlghEhT0RdMXuVrD2RxrortYOIj5jk1p3Bvyk0g
SaAJyIZGQjSWsQ5XDULYqlasnX5Kr2xEw6nYFBurvwLtUCDrQC+0jzsRF4MTPZorcVFyO8Rg9iTO
zqMSIEu1DJWzhlNfDHYaKtTLEbDq3NNfpMdkLy8LmOkap0ndXRo+YayfcZOcr/1K3s4NcIQRQBJA
AqhD4oauALafSis9/KRd+XdjUPNiEdU95SlFWTM/V9kFxQ6pB0/PAwVccEn78PjVtqOO6XuyCeTV
n530uGuva2CbuwBLdWU9vy/AZLa89ZEtWqZW8nLIuIuiYHUErmOXP0BYzqHoPQWurDL4URULsJJJ
kFyW9sLuFFHLgQzD+kYxN1qNoGNe5fovViLu/BtvQWOQh22MgM09hvQKzWOHcJK/3iBI78QEjcNu
K0jGzhaW8LCf5WeoEpMBt9rMFYzdGvhmARGYE67oeQt6ucuTZD/nJqCgajwZv6XmigarJqX+P9xB
OegIMB2SOLdhDMkAkHvLAlsG5UgFZoPjOKV7kMF/N8q3SsoFcCb398COdfBMjT2kiSC60HFyLE8I
Il2D/UTvchr5pl0BwO9SNRB49yp8jLRLb7rCadB5KxJw0xBE4w8pA+yYJc3yWYdiGgCBNJhzZCrV
ATPRtDbva/cCGj5ftIB2bz4+C3wDsoTDa3rNofO0U1E1p0fI5PHpOHKdMXC3vRAXQf52u56fYS43
6zwfpBCs7ur2zvB5/AVkY7h4g4IKi9ieqh9JSAlaUzVPxqMmJ2+4g7dY9k+0O7ZYbZZyLJhr0+Bc
mIWLUNkiBvYHsss/N+T26AzGQCMR2lGA6G3MZFPBDDC+6PFiG/dOpATGUPOFNGhHhwwZQyd9SLzA
tnX1DetlNrics6Mo7KSX81IHrikYN0/NgPvsVPpw9tajKWWRepXN8RxlbyhNmZ8A1PLBNutsQmLm
NESkBUE5ecoA/sCzVT/f8lHKuxTCQSaTfrlHXH16J0wy1PGh0ODVqbT8ptxKruq5AzuIHMPwJhDa
e5NG1mQxtXfSjZ96xD4mXUQoIrBQIllXPgJ9cbKgyOOVvfxDzKhRX7u0Qh+zBw1JziOgAISvWHQc
LoUXb4F9/azU4sBhUv3VKf/RzuKS1ObNkG/kEu8pfGOE+RImZpvgKWh2/Clbvif7vX0KuyHaMLHT
4M57m4irMTMeUADkTOJult5oSiYsSZ7LaXE35nrvV2R7M18ubHmF7sIRF39Tcm4bs/BqrPINVJcR
C9IH0jv1+WRgzbl5bpoksGaKVhdN8RrTSnbVOIG/r9liKRvqvIZylTw9lxjgaV4hshVl/OwZEwn0
3TdCbaLxXoTwlgGWOig2r1rVfnjJPlZVQl13SNmId7EswrxIUA6XrUeP2LFF2n7oiwNbdUu8DMK3
B4OnVXt0vGrVBhJQF6HZFja9lNmsTGJ8kriN8eLesaO0id6BLGaBb1tr1mcGhk/VwQug5mrC+yxu
tHSPvC1E5gm8MdnXGB1w+/YoqoPCe+lWxtSS1c2mCXU69EVewHnkjT5SXZDgKD/s9l3dgB1fo3cl
W212Pz2OeBlKLKintgfa9pPlXQUfEsZha2haCQTPEYiGkSBAc0sg+OXVSjAXW1Vd1OV4U+Lyx+04
aqTjLRojk0XX5NVpFHqnS3WgJWkEND0mUlk9FFWZJsvbtxhFQTbcEg40WBYt2AsDv9XLZ2r9Cb69
NmJBQaVzZ2aAONGDueh8gkWBDoh05BgH/rOgWHmPtPc9BVUVgoqY6J5/9/JDUOFi2lGGgv5jvyq0
0osQPUG17mAcFigo5r6WxsZEo7O7LJOU/cGM2Q7UGGxgGg846OamqsgqyeiqSAphZuDsAVw8+ujg
QPWeDEQEaiKm5KrOCIl4eQf1StJ5MqfRung1yOYn7BlU/RQHwcptYiQjBsiGW+b0T8aRD3lEhkEO
LkLD0FAOouGSYLlopiOksWgGGiWhrIIYGKLsogzfwbVZd6Ca0KqGzv6UNBZDjHbGhNwf64xZNM4K
lq4FJ8CKdQwh5CT1FA6/CtkrFbcKSN5BoNJCvI/f+ir9fYaKDXdrSlUA30Y+IhZB1e6VqzG7Ripa
Wz1cb7Srh11zSkUEp9PJI12LNSo+31Po+uV4cq0f433i29ARZWSfk49MMG61/5EA5mkbjoYJEvoC
+qjlV08qi+wNUhUeeBs9FOTTbQFcvjAkfgVp17we7G0+cOdSTHY1TYUs/SR/ImQRfZgk6rVyxMBd
LF84vPSu89gT5zTdy4OLTm8Il/ccAFHxciOcSsnuiBFYp8KumTG4MChWggYWCuxrDrN7HaOGg6ZO
KMaUHv4qumYyX9EiKZT2sWJ3HYKRtF5OtjBNpZ04/d/MNiV0dNk1lLTwdSxRw25tEpwKKfJodfmd
ALuM5MisksRB7url4Gu7tNyRmlzQffihtKFS/GDC/Y2bcrfiaonbT+dZPXgGPydlh6sNgJtx9a3M
+Osq0PozE1eqDlwu1RsFpACKwLgsZUeIEkx6rhVqyOJZXlCnAFRnXJXIBSAgIppxND46lmxqHA77
qLFwRiHngaKq5YVJ9mmkzJnLFfF2TeuTW7K7DhU3QRbmNuwTmtkudfee9z9AExXO4Pm09xSedJkJ
NIJ/qnxNTNbuOCSGvwcn8MPlgKLQ2lEa3eZj1sS5RSIrWZiTthSsDJvgjWDHsNDnfysTfwD2llra
wfs4NqiufkPljPpk4+WrIN9/aUX9Ufj4IPNr0XPPBCFjvhMbJEazMMvQR26VbNZ6zC6gTRcuqF4E
BgNVgNG3XhDqdUXG+GAR36F3j4v5njm2rnoIwEbOsdGnFham/tiX2zRUi1PSYLmDvaLMKY1kZXrs
3tw5Tt238UWGQ1sxVqhvC35Ahm7oglC2xtLipjwvjCDIcUMyDp3W71D/q7llYZw9FU7U/15LBoPU
c1dFn1aFRtDxRbiD2WBaXFvaR1YwTYSEnKGGIVk2FmZDk3T6Md+/500VYvkPzT3VUkJXHxqXhN4U
HEcFaB4yP2MIO0O4oDROPigHg6tYrLtiPL6M/HIbgD1G2NZcniDgv/K9l9rscX2ZYPr01aMkC+L4
umAwJvHolNO+GnD2JgTY22wtSqOveUZeueWZvIf+eBrkQu1fbgu2sTcsMROxZ/vS0rDpWo02xWwQ
wYMhiPzWkMkpkZIW1JTvG1crz97mgvWdnEv1bbgT5ZgCz0Jnm31Nq3e9OuJ9i+PVCYGch7Ko4le3
SG5fD4viJSlxUwJoedtSYvo9XqWv/ond2a08ljw4esED2uj0bTg70V6YGp5CVPsaBzj6xNxQxgPi
TG+1BxW59q1duVHeAQCjjb1CcARwoaAKoD3O/+XO8ccalmngNPGLn2gVyqb2/aqOXuH6PdeyzsLU
39FhrnjXyilEL4UrKn+y6bU3ff80nHgxG3Frol9vXTSSAXcou5/i1aFt0aDC09g/7sRLvLDaw51C
msXMR0EmIXv6DLD3oOSUTLs9HYRZO9ZPWDdY6nXQKMjHC+WgQh8a5bIfQO0bby6ov7hW7EBiKJUa
sDZPl8pIRF61ju8BTzDJO55WkaBYCGK8FKUjlT3H6NlDEe0pcf6pXBGaErkKsMF7aWbAOc0pQ3Xd
XofoKN1R1b/1B+q+lLOHr66UAwToYaQaRN7s8xGgqH4W7pcDzksJHHCZqLQCmmoN467ruDdzCG35
HXrNh0dslxSgDMYlgpNKqH2op9xTSrfZ+gyrupgbc7fPWtzNjQdQhgbNLxL1z0HqXV4qk+JTfaN7
Tpgfe0Tpx4rwbQpeUp0/+kE2+3aj4eyf7EN563e3uAAnGHNh+7ATsWJ+FD/xUjtoBVOK5A5kJkHW
IrOlZi5nmBM8tHBVw5GAQgTUyz/XCEsMRhZyGMwnCQbgcMCd6bOxmwxiJw2LoPyTggUbKrYLbReK
ETi2rOHme3tNq7Kgw1uZ0O7EFvmv9M+fFs0+VXDxtuqLQS5Y+pwgd3Ezy6PFICwgYl5De9/kQKJg
Q5qgqC5CE0MBQ6gzsU27qGbTbK6A2lWhltL8ullB01ajpSk8Jho2IXl58f1gN9tRruYsoBdBCjh7
p8U3Ki1wHokddl1A8655UaSP2nhg163UiY6A1+c3XBxh1bSOI6kZvULYklhFeh435Zk1Z5GwDW7Z
MMw5xDMxRf8XGnBlT0OGsM8/hCI+9XPyP4WZgIPt82I6B5kOhn/lZdZRjQHwe/5Bx9tEsgLLDuGE
1n4oLgCSd9HzVEi5KwjuTqgWTdv0hGAiFPe3Vw8h9Cc8PatGz/bjgJhXJm3Sq5oitD+SLIzyf65+
Ely8kzWKFFR3zqJiO+ftvBacq5bfX1dphcwWvVHY18ZaSvf2yRzZUBKMaRvLFDawZaWw/0Jvollu
yU9WUrOZJrxLZG3lgR+lLRzZJijdYT8MCoDVSvYdDnFK2SPn+FXWGXxMFSsKoz0wWTtj2q4k5WN+
SRopsuyGYrBrY94cD/CgW6Oy17thf1IBsaFYUtC5K1PrCKfUTbLz3dGZfEZszyXzl/lNvggLpoEu
T6vVcX5QbJ7Fx2PZyR/KN/SB9FMbhDF1aIfb/8wmxWEMkWjIAum7Z0ubuQEbykS4ghrmkkW7mH7N
IJ1jcy/5NebOs++TWkUDN6MAwvGWKL/CIffx+TolpTIXXYRnleg+w+AQ3zfCnwP6voBwhti/HzT9
3fxnEeirFDDGq3hKYdE3oTKIVosmmZVlqfcQlzbWSQT8i545hOFHizxMOp6GtTAWv4tos6X9pjUn
6I9mkzjgOQ1MfV4DVOzjkhD9ppJChi700t/Rhi49uppzC+zAR7wVB5OMixMkH6O90xcP/553PJxk
lv0h1l5Mvaq8dVamf49sMM2+tLEOQv/frv1pSHhfImDH2XeyPuoZDjKIhMjBLngqMZylKu/z79R1
0cnYSYhfsiNu8po/g+VGl64LfYS3XAMI7p7zL92xTpd/m1jxDreB3zVGdNYWk91QEgnEWcphCEr0
AuaTyO06e0SUv0t6d4V120K7is0RCbZrWFpquBtIP2iLUzmcymqBviEGur3rvi8Tj4+//4u3qWwM
XvROnCWVXZ9Ne04W9LfAi/pv5AASbGZQXANNt8Od3t6XbunN90eHYgXltFVuUGU4uAom0UY/t0uC
hnY5X43fsUjInMgSgpp+rFj9aMPb+7gLGS6RoGI/ErVN0HNaX/xhV2SAytl89pcWTnKRxT78F0qs
0xxKPw/yGRkBmx/YrgE0bokdEgqsxfYX5A0Y5WMzgFi3bUfmjkpOU6kyzvGck+D8ddG89oT8ei3C
5/DgUUKQzNdu9ZNBq1nuoyIpP9tIczbLfXcteCzJedOL+BBra2XyvHvjsjuDH2UHfm6kaByGYsj4
pmKHCflFlD0DAk9HKlv4/oBabV7ciRv70/qt5fw7DwMLW/mfkzDQ1bOc5s+72WLo8frIRZHN7Rn3
zyxSlICqLpD6PFEm/7HhaujB10Xj/Twtf0sPfqpH/DBkywS1tOVRl2H/yUALIbBsrI5lRyLgsAxD
c2cx15Gk+jou/X7N8NitfobdP185K0vSVfQhiSAyli4n6H1L+eYxIcCaUGXuAyj/HOQTkJL7lKiG
Gi/DZ8acPev4E68sNmRCdHdWhqdH5Vr5++VVKCD5ggTt3YBj8nOY6FJiypHDH+p2+DXwrwtvbg9u
bgvJZ8D4F7dvSY14mQaJYsbzCS0izb5oubr762H/p1uNJUf83VbiZQSfakUvQb1Ac8dLwLiSxln9
FmOLiQUlC1zdmFSa4GPAipFMNOYfMC6KNxXywPhc7zBD+IqvTC4DKujBzZZvOaB4zaWnDQlpPkz2
MznPdbgRwQFuRP/H1CnEH/Q39rURq0jMbpaGIux12bz0Wd4PaCG+cScpLDyRbbfJgKtj2tydlInx
0xd73nX9jF0rWwuj4+DEuD9hsLO5nE8aDhFA7dcXVTT2KbDBR8NGO8v2r3GIH0xdnuecDBDfxe9d
CSdMMi2Yl9IYA80966wJGmyKjiN8+EMv+Ev6Se4lXPemDL/Mo+vgVsRp5NgnpXjZjNpVRLUDe8qS
nfpFiQz5KY/D93KdSoz3B1U2mr2/C8mggPDmRUhreM4JkjgIKEGyeFDXPU71046F5X764QX2EIsS
mr7xGyyDSYGZwBN05+/KynWflJcIhvNuF4k5w+Z+PFIfziwAVWw8gMHUaXQ7bNv7PER0tquvcKP2
J3k8vxjtm79qykyTljMgV/S7t/T4+HnodDnLrvbu2/tUfy59+l9xTLUrE+sK4rXFDEs3EQxgZPJM
g/m1764o7HFYNHkbd8p5B/bue0aSyMweX/vSu3TJTfebxxcvQkVaACJLYZItws79qIV545WcXEFG
sz57gWToJgAc6gIQOcQ+mMe2/KFNC5dKyidrMN96pQPMVAJR2PECJUQNTanuVbOFIRHPVAl+YMk6
u4xX7ejHQudbISxz8LgC2Jr5RWf6bEd758nLtXIkRMxwQhWNZYdrQ4bEoy8A7iuoZsabTOu2g6b8
oZFucYTapBQwA56opQfrlhbhSTlrQapQOKdI8P+0qqsnAK80ALkKwXNEDjIKJklxu9rpB1VWbbpo
VoSvjoz1lSgjOep66j9OpVmuFT9LstbdrkYTcnCqNCgkg8CA40APACmRc0SztFGFGABkTQVccARe
WDCeX7FBfEuQQWI1mOjCUPJZS0P9O3+7CNjquICSpHrMWgIa0feTlUtWON+kxjRkeLTTWUSozlk8
j2Dtaahv6O1pvGl6KwAoXaDtXbpTfg73LHBNK+KdE53ucwa7Wn1aUQ9P6EhfojM+lYH/bNzUIMR9
udVitaSxPLhEkjUQ+VQKQaRa7z9IpGhh0FQxvAjavz0GnAvSI4nQEFWRQb5ZCTTgKgvEt0YwR8/5
29XOoc5Gsjlkf6XoMzGoV9doIJeKsKAmVygTKrtUjlsYEieHM+JZl/CZEnhtXLs7kW7NWOe3Ue/Z
bgMPlj7e45Tk4A3zlWZ5/X8XHlcV+FFzbi46a9rIh1kXh2fnlr7N7KHpzMX3g710IUIuJkYXwa5w
QqNedo3IsRKFtd8+JOUeuTML6Dg9ewuz4NxzX3cbNyrYKiblW+r8L9qntgPF6zu61Low/Rzq0eoX
SRrNydi5YwaETMk+Y2OQeHu0g7QxJtSaRoL3t4uCinhJtrchA08Zr6fxDtV2xAyTwKOdPCXUzcgW
/Q5gZVKzx5vD4QwTNF6Hm1TYdtDv86T64KVRZRWfj0NTdFJbbl6AN8gfZrPgl73Puyx3hC5mV94p
C15Civ6s3RkrDA1zFs7wVILz2IukkP/Uelouiy3xsjHPBr7srOfOnEkZJRyB6uAdHkiho56cj953
11Oqa4eXs9sIW9XtYg30wndQskJ1Km83bjnvpBt0VzRWAcBmcq3aAb5YplCJnUwHHMNGIoSgI4Ns
Fgibad3Qfp2uLxAVB8Hmwb5gkgOS+YlEKE0V93QhyLkz8Sy7PyMIR7N6dq2mONipL8T3H1SjJ0U6
3MW5j4to0Fu8G4mNWI7Y80c7zMp1MXajoHcodfxnZCoCMs/zwHO+ImhGtM2Q6neHX31Z39KUP8i+
LdIbSDnBWgX0oeZf1raPmK6XQLABMZbiR9WSt+8cmoNW3/iUEgqHiaHi26NsjRD4meksLnb69R2X
O/e4o5J4hIvsgz30H9zkQ1Zd7A44Tr8xjCEIM32SbTFWOtnbKhUEKwRcFiJF/5tgJfqW4waV7lnn
gAkYHgN//WoID9J/BsMWDu/TAZPPipRVOyBv2Uj5Ja7fSzokf9T8ukcKClmRwOj+4oJEk0dqz1yL
4PxFGynJQiIqj9BXavhjTqhHYi9rCwfklarxxHiQ80aphkPUNPTD3ClCDDUQQgYj/DoQwKLAKaPB
71+sSAUDQQ+k646tIMjgXIwQEVs6NZSdFpo3uFHpWunlYt8/X9arXk/OOloyhsWgJyE5iX4Hn7bt
Jcp8JddHNd+07n3JA5THddaPqamHyISpZP5jvkdMW8KOOy2iy0M+5aqv78TZYdfd7dN/2yWP1wNx
5+j+Mju08SBS/cHRIHZ24B+4naHlB81RGzXqZyxPH1uO1gP4OmKgr3Hgdh0ckR7BsnVgdudgbdw6
nV1zJlq0Ufhb7rbw5cBRqhrAI5wFIEeVudSzHEzOYiJ7PVGkm01Pyo8FYX87avEI/DZbUy9ouS/m
htYmjn6C6kKX0iJr7yW3otBwGXM+IAY7AzvR254YPhAqBmdjD0BSM+ImZfxIDs/fTkhrfNy7YQxk
OfowpGv67nI8tFTlGCG9pjbhon5qPCvR0gVKfFKfS+FqBhBIcDcDYEXI4BTlGyyZRd89c0Z2/aUT
Vw1gIIzB7/NARW04GjDt1IejcpN4tzrufVDrx1FIj4m/BiFY7RPC4HO3eAE9LkkSB8Z4/YG15kF/
9DwqtuFXVeo223nulmog76tW0D29S4HwzV/4tc8H2/Pm1Ro/LCF67sErNEzI9oPlRwPS8hZFbi46
uTbPTW5ghdpoPv9tHxDE+GcBsntiDEDE+w71Q5CTDbaFGSHuW9yvHomXGJp+qRWkW4NST+xwPenU
XWTVA4INt+BUoF7L6hXfvyEXipZ2sIyZc24PAIhyo5bS0M7eaIpDhPJpnFi1fqKo9kMrXd8vCyiI
DtQSTvpgYKvZE1sxVRZGWN8+qn5kTXcv6heYnY1FVwjy3y2O2M6w0AZZv2NSigGWZ/muGy2h6nwY
EcacQYTYEjDvaG+EOjRtXZ5Z5vgMJyRB2OnIWDpIYL8ePoMu4ITZJn3PBdTRfY8pnl0eCs8Nh68t
iiEr7qvgC7sk77hCgyh6RyYf9MZcS4TeA56UKl8px/PBWt72tPEKHYzyL0ggRe+MQx6r4tD2fekk
H/e3D9tG9iSAgAL3UUYQE7f+4HCIkGGbIpVmfOhkfKwqTWm8oxLl45fiUl94F07R90EWpz6MDDm7
EDjxuGA3pfADI384J1WpiTo2wEqBSFGVb5xYlwsD3j3cZYFK2PC+NDumt4nWJsfCnPQbTiFco2x+
6g34sNK9IY5oaI+r0Ts/oPCI1E6oEnChmvVqp+wSzxQ9b5lEdXGfjgg7oVrenObxONN9jB5RqEfA
GgzUOEnDtf5FQ2wPAh53fv3X9/RcTQmKr+Ufaoc9DsC5Ia7JL1Mh1pfbKdEtgGoClIpTHDcI3dtw
TC8+onC/Kz15zAhfu1bTBEiSa6JizPe4JknfrsZSOzu3OH58GDJwNx68cFFln7bok+rEte4a4/w5
UIShxSgtDLBJlDhixPiYV9M7I5oXrj3jJCU3qQSwSosj/zgijU6tdBxuczUcq/9U2ubAVjtiI+lt
ucMqWJGaix1AHyiqBqeJuEcMWmze3otClX0vd8o26YeYdXoYHcifY1Fzy1DK3KZYzuMCr4+FvrqO
uqFH3hm/5R/LWNUzHMdZnBWZHm5Knl8quDY7vWvZcRjUPjTkOR4Sl39PQtqagXGXBp1LJ5S1aLiH
nI6bkR/CPcGvnGyTFulgxvl4skiCSVWP/+uG54a568zDLmnuC9fm1I+NH66GaBOVm31AXwCdKR09
HHGcEAw+1Ljld0Sq8Y+b7PV9o+O7jbU9/TSExjHG5tUPGMZdGjUIMt8fiIkx4+pmWthvlUTs59yC
ByhPn8kLEVSWeNRY3aYKLvXDvxW0/rgYUzRtc7JdKoBKjogoHatCMuaC8tID/NW1aOoIXatPxfu7
PdtTHOQAgwJsV0ee5NuTjxjmc48PAD4ygmlg2s4fjz632ce9TYQSakPmoIl1HlkJURGu0XoWjLk+
sSoK4fdariA8/pH3TsRlw44aPKCiqqkci0ljlts8kFYq3aQHOHKlJt+kBru1+fvLzu1+vzUQ7s5g
0WfgyL80TdXZoHhY5qSbX35RNMipy6vQa+PY1MhP8WbjaJdyo0wuZXsSd35B95WNB3SHgy+4LCCB
8uuXdd6hnlqJtpEJPUlQYYUvOrgcLhAHTZSnyOaCJTc8easkOM1eHXLx5FF3hTdk5FDoA+c2E9rx
sHXcOQUShFRwQ2aEil77OzfDS7rKjQJZybKWKOaceW/+Qv2TcBUeH6ET9uvfZbLlteStTwgOk6/u
ahKO9rmQB+Dqy02FmNRl/vJrZvbjNWL+bY6KiofD6L/uuw84VR1kCUIWOwV2RBE41huzmz2zilCd
Sz5gve8ywcolR1rzcCcJU04vZR8647Wb36E7YUkRSVYBmdKOIw0Mppe7cx93dPi4X3OZpTzn0CgH
oJansGLD8tzNNynt6FjFFgOcqRvAkbWGoEwUBroD+FXSLH8doicmQpvRJs6ixAUF+turOWBU9jTO
IOrssu2QVpYTIRvtkMdzoYZLgYu3syrqvLC/DfV6eJUELeyk4gC30DIK0lNARLrEB8yYg3Qw1WbL
u2AjMzSgLcMSu2UInOpKF2B0af2GsgiNxN0u5evnqzUw6JRwtuokZluDYv/A1aYLNmTQHqPLg6DB
2R/klzUguOf3ePHyT+ujMEcODB1YRMxVtFgyVdyH6UeGUMdMH2TelWHjTKn0AWjQn5Wvz/n06Mhm
exyvfXc5DrbbXuzfj7TbIDZQuhNtRTlK6nx5nYJz3ad6oz5vqR8luCrru37jSZdmSWAXFxFr1tlW
8yrGtaRMKSFXe5xNyD7RwE0l87Gp/+vhou9H4rmdRhJ/emh7R7tFIAO9mPWe9AXivAEPvpVfWhK5
DhploE5BrYPx3SfbYIvj5vuHeAIpQ1UtK2UTrg6ENmbz5qwGXBlDDHfk0AWEyzwLdtn3cv1vkn+r
F8yaO/yZYfAk/HeiJmckAFhMJzkitlS+bf9MDqDeVPeh0xWMQl6YVX7iv3E5jAzu0uA+r38o0jeI
qFC/r5vM11hzpv4Xzvt/P1G1ZWcp6mjt74tXnRCS9vLzmqxEOoGz9ppVq4RUwDwf4ivsg3nA5bXR
csxMWYHPtmTHXEeJKNCUIH0Ax7yUvM2ZhrDcaQld470K/IkzXxwEv7kf2Rhy8sZW83p9eSV9mJfF
15w5VKxpkc67LrmOfYCSchueJ1t50BpVwgoBpN4FF7C4Yir09u1pwZcKHYN9/5Y4OPXWKK6uttwU
0VFrHBz8hsQkG46sxFLE1xh6LsEi8RLKENawiuKUC3WiWl5ju19QJjDha1MqYswBs6oMpUF79Vzd
EphvhY1/rsvmInsTpyAd8ZEsdtzDv+HifIEjhCWXQa8pg03aBSqHdbZhQ8svT7WFFxne+c6r1Xpl
qkmG4wssiulREtguFbCUl9o3PoZJjJuTxxxf/a5ZlKpQ3Y6puXY9E/xHOP70tuFco2kLBlIWinC3
HwMm76MSdO7x8S+r3lg92N6bXXkXKKFOfAUUUrs+2jeev8m5zCepEjxs40GrCY6bx9b2chYaPsMy
xu13WxzX3V1mncxV1bunysMgyr0zWWSkGJcsNUzEragWGVPvOCiLXCPfkgFxDgsjR+sBypoVCwSX
Eef5/ypmdwNzSNVHeKQxXa+Lm7WstkqoR8A2mGsJw9t3dLsMA66gYN4DI/gAKLOEA0uMGtdeXtHG
fEqIYi7lr4/otViay0ouLnvhRUza4e3hJaeYvviHyidYOzjK3vUdMxfCJWN8dxkfIIHGLxIq+9nJ
ju1W1fpVRy1jWGT8IycguMz+FGB+zT8fmiC2GcKIolRlOnMFAawmv8zHg2KN3CBGHtOnpDAneTFA
XRzwcacB1ije6OIxW2e9BT/QrrMuvGc62+nps7zmBcOts2tVGUYTOQbeQFfET1IKFn7ptzoq69kN
Ss1TYtbl89ZOo0Xhut9iCv7OHZzFvgkSTUX89uIc3qRBqbpoBgAlnBrXhE5yUabMSps6ZpUsFdeK
JytXYARRle5zn3MV4x273iHyhkX5J9oWxDGOBNba+er8BmiJSv1dDpTUmtAYys5efBgkX2Iakho4
0YibgPRGhCcA0f7T2g6C6OI6V8Wxo1Bk9BLcanAGI4gbXz6S3U1Uq4rT7g5+v7WdR0sbXBJniQKf
y1L2eU27t1J05DWeDk5r0+G+UFreu2mtWswm+l3m8YpztnQL7+7UZ4p26TXV+l8W1sC4m3ktj1KX
cA1UagwR0D7Bh/RWQw42Vl3ULzOxhZSUCZC8mxL4i0TawzOaOl0rMzgtLueC+iX6/Xb8sQJoIDTr
K2i3ZgpwFHZKXEJedSI7WUpBvtY+tnpa+EwtSWVyq8vSLZq/zQBBXyEkqF2nsIcBA/peZNNZK4BP
qTeRxCrMQEz2zQT9ulK/uCx1szrjnBHO3/e8mSvXow8nvXRVYlNAGLWplag5vid0gITsKPAl+8UE
aywLplrx1Le3P8uHqDaD3WhfwIDqJzzn6MUt74eUC0jBrMN3sL0ClYUcMVF0Jmn+MrPf1lGjtxmu
9WhHO+YQeG9Jswxhk7MLjXdTj/r6cPhyUgxcOvd+8VC3iRHQkhLEyPqglVT7P/xAsym7wqt2VkEX
frOC9UtJm+CoFfWS+hUg2RMcdr5jJz1WtYnGdJvfbPfaJYQddz06UNf3SPqT/7hWXKMfV5zCp4um
0xpE6Fuog/5x4be//5zWqpSFIk1244UXpHaGAi6oErVBQP4azyew8YZh67x2yaakRYq8GpuHfsCm
So9lTt75duZoDO7lYd8b/AfCaLhtWDdTUCC34txHoUIo+3CtcNdIhyXqd/SJ5QroHnuXoS+rqtzg
yRsnJ6M8b6z2uHFHAres+TULJlIYW+TgLttcyBh1PxA/h29BFdJGwwBJ9mobk7WKPGI8Ds3U3Sr6
Xy7M0/AylZ2m79IG6MIpEhBszYu//a6aoe/BZO5aH63GWW9j5B32fWSRYVPoYO0UkRPx71Asfkqx
Vzfi1ZXyE+IuummbOEaySzDQJzz8QxsaJktbFHA+/rZ58f3oW6ciGiBT3/6NGTDndsb1zhjuc44Q
xHprBN072hkUXFXLWLDOJomjVezseSm1kUWmOvy7KpubqtxqYLKlITiz/6j9jyQgCMEXemNBsteI
8ApYUGHsTM/izdYs6EWHkLVJL+Mb7IKC1zMGIhZtJfXGYkqBCRDj8uplgOgh92saagQX8KamUCVC
3hM/KKv2Zx5gzbSp5yuPDZ+CNOmF9AN2QkxYCSV5JPHGysXtAg3TKD5PIkh9PbWYb+AyqKiGJoXc
4nQcDkQziMz40Zq8capywcZwjP+2sOh1AhD3sS6+kaxkU2V8LUDxAOk7zhnBtdeb6DoKAnO3JXqt
rOvNaCo7IIl6QWfvDkhaNbQnNWsw2orzZ0CeZb40dGRo3E3Jm++6/AL9pweq5a4gTHWAVcn65cqR
GfUFS52hbD37M9YKcws521XakDXmuyizF/fibZ0ohWV0GTD1OpgckW1lg1EUQT+dIM2qgEKqu3mk
tPNzwWy6g+JFSKWw9DBN2MPGIk1IrwU4NIx913nXdCSMxyyH2NkiOavMoJ5ihqjqChvfFwjyfgMg
MY/gpiyWgEsoGxmvALueTuUjYxEQeIBw/qbtAMGhLRGIJukmkxCCmzdE82l/f0Dkz0dqMWz/M4cs
lv9sQS3YKErdcHqyE9BoSTDwPeLrA3coH+GOetP2o+lpSuFCwsFU+DkPsMK0vLFUF5SKmQoAJ3tB
SKmYm8Ypad+2txpeMIYFhQJcWHP+WUzcBlScdtqORzswVUctIJYOyXTPNHBVOciCGObGC6qQxR6d
WKnLYQ78NcoN6s9fs8vDohbI3SVHN4XN+v7dIypZE2cRmkbefJq3D5u4+Qb5eY1lQP2PqufSB0/m
bRu4yspIcr6ZfYn1ex41LzPySiSddrqVfTGThfzAeo/HSANlrz66ag8VnI7A0exY7L+HHGR6JV8s
fOLBXMdf+MN2OuynxWVUDaXCpRypT338saqznNsuqINeDIdbhFaeKIdJYshXJUMzF1vhaEeAIise
1gZ4JOXMOomV8lAzpTOPasbY+rqHFpgirWOahzfvxkSo5eu1dN/KXkx0SQNv6LukqvLNp6kDmfZL
LrwNdiHr8ZiJIvaPgxNM8308ozamOy0Jz4UrqqVXp4R2XR238Bh/qnQ1xt5WCiJqI8n70FdoHY9G
WkaxXkCcMhYUiPl3ucndUp6pxi2UB/Hq0HF0F6e0o4uRpleFqefoLymtU8w69/oP/GofZ9uSJ4zu
MipRHv79LuAN7q0BfjXAJAc1YArVnQxe29UL7CRhmrhS0OhXpoKBk3i7uWVjTGuKHKvm/Fw/uC+I
qxnD0QrYrj0nk/2lNwX+pM7fvoivz06t7bH14Ln0BxpzL+6ZNDdtQsXGc4mtS2lkh7qBi5rP5lHl
SrobX+GgrrpKzLS8i33OKbo0sIAcdZFpBWZTb+VcZK37iDgkKk5xjS5kwtz/hV/DGaGR4+sGZyCj
0r4nryTlAwRPRO+jVu2ShpIXFxzrlufYtqu+9OUiG9YY8/ZfQbXiL80l0e1X0qg8QFCX8k5fMwYt
Zjfb+3sjRbh5O7E3CvXogQaTlbPsl/KDs+HYx+j+SpDijXMoEcRsXMTTRrl/Ur0VfUCa9hVkeYrm
oiJFGKi4nvfFslQ72/MWlqznroMjSsZDA0Fb3Tv+6PmXu4KT62nOncGhoNjyEz8wiFVQCXnxbnXo
HSC2OTGc3MDcMFX9IWl8hg/wyAnIZhx6LR+vSWGTjOniRKZl0JeY+CHJ8PAsEvSyaHGIZXjMSuZ7
2YlBohHpe7CZ2kOGI0UTyCzcCwOTVBOMzLEcL8o7arwEgKLJdIOLo4nvOqqKI+Xk8251hdkuXp/I
HDp4l+X/CspjZHyDO9g4gBR9osxJ6/4u9cu6BAoeaO2wlMIk6UrmqevZZsxHu6Ri/M1CXJIEROhm
iJQIZQ3oCK83GgZvUA2cl9ytN1O6IuxWRmP5tVMjjzWDb2EXlQB8attx7B1JCV6qQJmzfN7pNb1X
T15e2HZI+RcfKUDWtNoOHGcXWUSfWDCguy7+OaC3+Ec1Odr3LRPxZxYCPpvt/Bp81f/rptP6VCNO
TIu/fCe8ZZVKDxeeWkdOlWQDN7PeJbf79g9iEYsX1GKOSDIBprvSBpYAR6f2AXulIgxp7PCbVMSc
4Q/vR01set8hTSaMxwfrB7XAxphJds8wMZ9nzgYk3vQz7QQTGLQio8z079w7rh9gTrVcTIs8evml
u2wiYIEx9gGMUM9BNy5InUfAGlwTaJIcBK3qmXbg792jWXfL1x9JxR0vtMOIh7ypLurvg/X6UDbx
PgC+TgLX1RwuUaSXHYAJqRA4ni79d4O1LNGgl2ZmlGo8+Ej0WzqTHln0jnWIZQYHjPRzPCZB5ox5
tyGf3M+UsF0rJqgBUP9QiZ1NIRTjJcnckLvDzGYt5+On8GqnXxopVaMQoIfI8lj0rahcT/kCvBm/
Pgux+ThheA9eqlIIUc8e9DXb/7OIHUFw7V+3b8zeD6HaQ8biEbuUw3qXtm7fddg/B9GZwMNPfbVb
ffjss50VxMW52D3azDkcWlfZ/opxJoQeDyEGadcTp0UYqmp4y9poDHpHaY2dkpSfKWf5ljqVYSCn
GFCidgYYVUCNoopx//JQa14w+tKBGRzCTF1S/Y/h1JkdPJZqt8E9SBlcNsMQLWt1N4ZEOO2N4yyP
OWu+12KQpHHwCT3XEspqPNVKQb1E3AahLvzA1/mnFnUDQJcegBzfV3zMF1onq70oF1qZ/khCKiG5
IX2T9tUR8ltlWb5R8Qkv8ab+eMcJxQ7b+5TnbHQ/Q2BB03vSyiLEkQb8cvi3mDEr8JhP0i9VUA9h
jEJ4Y0qQ2u3Rj/VcKWRGTavvDLoiynB2JeEKQX9Fz8OyL3Hxbny8JN2pYeHQRv9X76Yr3LyITk03
7fx9IqNCwi+w7/pzw7LU7Rf/8+JuahLdfv0vVTDepQftU9LzNxvaW7I48FamHIn4Hu0wbRepekKg
huYveRTQAO1yBeJM0t+vTt2BCmY0hsGnJrtGR4zTJVmXkq/emoMPrHRIHIsXF104/zQ57MnmurHc
9R/uqqsZIy2exicRqwscwnibte1WbeT8aBoC/vFgYZxHqtYJmwAUCMNMJJCN+CSIMlzmrq7weAvd
1u7lxmmXdnFOrNxYeWIcGu3VEEPBCA6KGYPVQCvhfsGgRq9G6xvFH0xYRMmUJN4Ux9YaOU09ER+B
aTYUnBP6UmaZBFZMIJCGR2TF2KnbbIojzurQqlkft1wEK7TtAS2ovrmyNDUuumpK2T0SGPJGqFH+
QEcr5WfFL1LP3CtOlLLqoxa3YuIi2NzfFLsRRRGbBXAVMFo0ADKhzKbKRQBIPSL1e7xHUVaqfFbP
wZ+gCimKbMVndEkIzkratD+QDd5QBI/7EvBIm3SpDjh5N2h03lGUSeAl7NfEIj1qDYdr5EktgAOX
u+B12Yz5axyEZPLzVzGXWTGmwhMzng+GHdJlZjDqpWLWZvolV8uVxGhUw9OcF87BA5SN1udNHXfu
P2/CuOJTMy8MWT2SbnMIzWsMNWGkJ7V+7D9zfilw6VI8TRR5efyLBjn9NbC7gBnavUDPqnxQ/7W8
JIQlK4kOrCDrC3mo1ffwuJ8UWZ2Uyq8kjxSPkc4IBIwrVFnYtutCiTnf423LyUfyQ6WSYBqz0cm0
5mLc1sUnrEUtKA7MNtaT3Iwy3z99yDaNunM32z6mnZ0mRVNG7CannPgKdwKFrnyIcEaowqRpjrfX
qBxUP8aOjNjdIe7zwaL91bxgVMWFk2WVQQdOOm6Mla2WSKd+4xoj/QguAW2KPRwC5Q2lqDdjZQkN
ETBHsH0CnAxbhu12lkrV334/wkSNVAoZ6YbmUSYrh2vwpugAVuSmUW2vl0VhFo9FOxBPND7/Jb+u
5N9qf6Uw1dfTqOES+FSm1NzHkiKdB+KpM3ctDXIbiiik21pBaj4Q89PXYm2uoLlsxssEe/4+xhzz
kp3otqTR+7ck8FqSmgx9zXw5J76h1/j2o4WcQLXfWpqCc9gUbNI30kEVybyeT5tPHcrppBUHsxJf
pNvjdtHXpp23J9Z3xIDzCbR9K6SrLcnqtsRbGwaAeuvplEkO3s5Cj7cf/JsosEtzmaSHgOVv9qQq
L2crZwKaubJUSIo4GKtEH1bwU9+u9ad1Cr+rlla92YUBreDy655KO+HQbEkEkb4xYSfX3nLACmPB
v+Bb73QaHlwNDpato7DNQ4aT+I8088YFJA+QEGW6Ge2fBtiN3ag3xv7iSGppj1c6QffPJ0qKti8z
vDdV4nPPsL/gRzU7u+1cBPtG3V7t4S3kWaNgML39Q3gkZyvFBVESeBWNODVDj4q5Ykok+7i7DlBP
yg0qvgRr6FYZYZVjOj1NGSUP5UXHU1mxeMcAP36QeujfUOfSs2HiQa/Df9JM5jaSVrgJsHci0SS2
/V/tzsubvdma323bCM7zP+JCvZUSLDpNdabRG0ltfHv8j8FTeSR0YMaZZVcuxO3uCrdsBPSVMfdc
TmJtDhK3u3qPG1w7PBPjdsZfcZ0m0rYPl/zwZm9jhgsEsGTKIdjzHldXj8wc0EzvZOLeGhixe+yS
6u08/FMPh1ejk48lw5DCW1c0J8aYyWp1eMfgDzaK7V7S33cn0XKdXowtoaY78iZcpxoucqI34rw+
aG90tdlTxxeU4PRZzFs7b16yz6qexpOhJ+DES4hGmEQv+8FlZN+2wZYHhl7VKR8lJED3pda7mj1/
bVflWaCnytE7ws5PVp2fLMnWfKm+3tc8aRzZFQsCiNEBtlEYKSE5PDESIuI2JpX6BFqpMpBAq3Gl
gF1J4ULGRBVVvq+qgDTvEIz0V3LSrXbRUBYuaX86o5FqlpqeCfbCr9uGPTDs/JSkS4vH6/nNTOXR
+TB0T6HH8EOKf16yCh8QqwYPIekH6foEMP7E18I/DQKPP97hn4f5LAHwKx5m69Y25UMgsiRI5/5F
mQ3Xn5niE7YkPT+LmQRJ9tlAEy84L6dKerzjlAkDlVzLwaykZTP9bkFNSIkrYoW/XAd2ZXzV+4Wo
QOFY9BRtXmBSfZkPMmYUMbM9SFW9GsNirSEdGpVMUPqOYXLrMsXqUhmHdbcgGXQArlV0lPhNBcPH
jkZAwLpbzRBNUfsOzr1pAT18/wWzQNf5oX3In7VRMJZZMA/uVV5Kb09iUZxF2TuNdxqzGeBuOHKC
pA/6unJDvNu+/nSJxDO4j1eGq1v0/MGssyvHtit9Kl4HOP4gRxqaTveR7EY+1cOBv8AcsEm3T0kv
96ZRHdE7TIH+hPUdYm3l5wiaLD3yy27u6w2SaXPXiPzXdTk2hsGN1ntdsxictaQplfXkdZyheEXI
OSvVzoQckYJt6fDp467KPeGdjIuY3TndQd26JvKXgcgNSBOPnxfOeQRe/hxrF8mD1Sc7PsuAB/ig
RBIX+IvP8eUqi6l/dgJvfbVuGg/FlrJrWC/A5IUN5YVVqM9UMV+kpwdjLyGRJyrWV/6sBs4iwTYn
kxnFl6SKF3vmS9V+dLj6SLhf+cuLiJ9O4S9wwRsvXOVMyCKL1JFHQfASVu3bPBxriJua2Ew3Ro3Z
wXCGd6CT+Pmk69WWZjOoN6osX+ifu8a5F8HCNESqTx7Iil0nY09DMczN52naVRuaR4yPYGMPmnq4
GJfYW7H30ADRoLeSTGP1qSQg0tV238hspJRwJ2hb9BdY0hR+vSHrIp3pZjotP5kMo3sD1W6B64bO
ndgJRJWL+I2+NIFNrCUlovWd9TlLRmwWPWPbpmpiQazXOI3aePez7hZDcDocGb3jM05iUjQNiTgL
XXpRompPq6Jkf9Y3NIsOsjFN+c8WLaedyr7NYFkpDcNQiPbJnM6nzZrjIlC+hVE7DmrgIczAKGi7
GV35cGDWinsQBUqgvSf3p6xiw4rIC364yo0l+oneizAy87S37o3/LMdrqkmRMLUsTEpPvSL1lUgH
oaluVO1maLiZur1H49aNIuvgwBYytY09F3uva6lEBuff0ZXtiJFoHjNu/1SkxnI005/NbBroQ/ne
SjOBLGArkDSYjZNw33EBocXJ2QBZ8HVij+GeBRiMPRQxArKLap42B/2+0YMBG7MzYGj/T47igJQO
Ez7hihsL+/52yYqrhqW80PrGuZguYOH7WA/k5jg7yKiBXAKo5fbu8wPngoM33Vhg60wzSoVlu5ik
Z5uIWp85IOUtYFvTJ8Y7yPBjDYEXYGcozlV0eIQlMo1qXbt5R+lXx96DYF5CYCRlqNMOfXgFkh/6
71rBBhZDscFHT/TjogLl9HpSJBwiX/ux6YD0f7G5U2apV6p6zt49EkoU8Wr8k8pTdc/8vpm4MufH
aGVaS6JZ/04k+42thpkruqlTlDcN0V1aMW5cpy8xtZUjXbnp02XcwRAqRaZNKhaAk4wEoLkutfOX
SgPvcurvuFQoWMT/0HNWdWk4xvVEtoOdzMJD2PHixXP7UmXP18fGOGFNSDH7jkiCFbDlfCqr6pTP
g4TlQBTdFJznTg+rBQQDWnmUPIXXOBkKBjCZahPBdzDdX4Z7u2WlKMFU3KbG6fCC4SK3RaiE3TVn
rQaGSwgp3XLW/Ocrw0Pg0cQFmqqH0tJH0J9PzQaZywH7izRgbz20hzMxrd1LmRfG5iGvoiizAM9c
p9xNAeMnWCEKVakJSdM0rvjiz+AAtq2juHY1Q35yWRaCgw4QEowhN50zaWcxGwWePYBJpmRpVGZ1
qUD38ap1Do0kg5XfFrmDNTctPf+zsD2vVDbzpb0QZp0puVVji6gNLbq29pIUQoPicfLHPjB/GLf1
4UHjy+AeMHNsNlTKGEAVSiaTVQOIU/r62kcFWcGg8Ez2QMuKdyq6lEejdmH13AtxDDjozNPu/tFP
4IsDKDS87SSPfr4juMYlNjdiS6UYchs3EfqEZDJcxjuLuKv6eFU5aTaM8EGLtKhMXzJX5lCWbapg
PPvhI0LAcSTDHCLD7IQhdRr5g5i9aveCOQ8Yi6jwbuBFPLO6+TbZgkkOsn7EdCryBYQkIV/H+9Gs
uPs+ASyQkSJt1qDVWxCU1trShpO2D28zZC7vULKN1MopTuKSFFuiqimjW26lAPZwdOIq6WDAcBOS
RqDBH6Po31V4pwgZxACZ2sHtjkX8LPOWlygBKj7bcRzkpzwdLKfFAEaOobJwYeRR3SvVAj/j6o0x
yiRbVCuosTARzF462g49/Vjd4XkK+o/mEjcPKuj/BDxj7kyPtXdfw/aASR6ueKPK9SIWw0hc3SbD
lddVB7eZHVrIzmT9jyLhgTrFxW1D+87wMeqNfvAEn/N1YJyp8fC8CJEkWyEV44IBrlfDszsfiRfs
kPlxpFIROtYY5lIcg4tsPkq/ukGA3TlAEBB/9T3PjcsNk3MIyC21yFPvsSGQ5FCABkLWj+k+tM+9
ycOm2G5Wf8wRACYP2kqn862q23ubvepBbFOua6vubFLpqXrtayfPc3w/ocDKyDvUdOo/HRJ4eAs5
eFkFLscys7/ZcgB0vZWT3W32wADr5L5h/vj/bG2RZ41LOr5yUF9N54j68DG1Ajayn+WxBsgkMofZ
9wKbU1Y4aJRwQeiGuzSPrufPHHsLEHCQ+pdjGsb/u7Qq2im3or7xz0hWPbYEN28GLefFiAkd1hp8
aqGdQOrBeCxLM2YmoeN3G3tSmEd2M3oy2TUlzntTB0/d253WmnOwp42FOIaxTjlTp6bo45tYAjE2
iF2N4Cut5w5vl84BADk2Qxi/z1PuyL33/h/m9uNSQQj8layG1gF2bZJjXkSGfahKP5n22uSiP7TP
nC+xoSp9dwgm/sVxRKA5VrMHHhGFh/IiEMhXI5tGHxK3oiWkBGRlfOxsvWNhv0lKmAkEyWH3wmFy
yp9EpgEbhQWH62bAXDlVx8qktcVDOptX2VMBFgU3yw0A3S+cMoRTnJxiGdOm9Gth+RFLh+h7gmI+
y52EFPA8C814OKSsx5RvEHvu2snE9gCb7RTgPp8HXDyxwbdS2bEz9gQJTgZKbSHm5ctDy2vXTOtI
HxrhTwJasVWF91awTNcBE9VpgbuiOz+nEI08nGV9SBevCB4Lkhn4wlSDAQupta+Z9WEi+S+egsbu
juJTwg3ybSJm3egmLDQriGyRdm+gKE2FOX/K9NWSQ4QVpTAUYdtZkROQmYXbpVSlXxKf/9PfNaNl
N4Zk9KgaNrJegSM8riEMPL3p0PyHlmVhRRY1Z7RxXoA6AgH64NImU+/rPP68Xr9Sk9/v/RhIVXbT
f50Q/cpxJ8Rq6QaqtXjyxa5AbfHn51vAPWu3Y9m3x0la84otVfXw7//fU5Xgy0yjQHT2RfYNJNJZ
UJMnKVmoxFqfnjjBk4flVP5f4WOCuvJZJb8lIicGt4oQxCaM9KYTtnFntn4x2PK8dyn39DiRUg88
X5ydlklvsMs6HWIju6yAleTQ5Z6gihKEUK20lzeFeqm3AghZMffZ7FRs0pcWwx5W7IJeKeCTP6V/
2EQJ0Qyoo0r2DYlvNatXyP0oqKcIsiLZVPO3ljbpKA88gZ69iRTAuyU5hNJDEXEDtqLrRUx6IQFd
ieRihhWQFwY5Txht3noy7ShLwSfKO5zCdyMgoSoy7o2eLopCHuwWMpa+HGmwTkgJW2TfxGvtRbO2
VYrZOJOARnX0zf0lwo+zjMYtgasYoqvjtHALh23GRiSmPh1WfJvnU3840kdRA1kR1QVUzkYYreec
RfsJaa3UwalvJTbGxt6hUy8bVoG+NievT4ri2FZAxQqJmS55Tu/Ue8EmOsAEQ8qaw+3QHf3w08Uo
XJTQ9WKV60PLzl/L6K3/gKD809QGku2+vkUTffoHHQlzt3W2w+IPOc2TnHraQCRWnzGB39v90LWG
e87VL9AECmrGId8zEhTIr+xHMqRNFoESR902sxL9fQ4beFO1pQ5tU2F+/zCYWJbbgIim68jEPd+4
7Zssexr4NqdoLcRlG7Gqk8YyhbO732I0kgYKgAJxVLyD/mTgr4ASd6yS68yL4d57OXYccmBbxL5l
HR/Q9khSasnD/ZtBpadSJDmjdzIzJ5xpayy3JUvC30wGiC3N3V/YnpOWSdZRTqNpsNtVZhWzUukr
nvuUmKxZxnFYW1DPI0BQb5hxJO1dLznlWJP1kEyDMmB47bLTS3I4/LwZDuzC9w0eY4z1Ry6t798K
EmIl4DqwNAwqBTypapU1iABbzpIa2DQGjT+m7dFO67U4Y+WCoc3cYceT/J5/WTeQjDmyfvNQNgte
7+BMO0fmOYDEYkIidakLj9cHNIFjPH1LtIjoZKhpuH/jMzwgy9WdLYedVXDYeHCsvT1ZOX5v/RyE
dj+F8Cbn2pa4oS6nIKnT3jchIidEYkQr78PmsnHoKfuSIdV7biz784h+ojl1dab5ms6w7k96z1y8
0WFdKc+JPIcqDliVlNnvEXlOUCtmhy8gOio7qjrzpZHOoQOTwbftqHy0GUZXmsliqe2ZIs0uW6pG
ljdubqtnaaMd6eljGa52vgwPfkmYZkqfK3N3qtzPbHzh5YhiVC7kzhsXzAn8DB5sbl1caCc2/jtW
ofl1bg7z1/HNOBKYGKgyl0n9YAAkqRvsGRPrencIJSfLDMkEp3O/T5ORJdX5BJ7B4EnB80TpS61F
SSTsQWjP8AzfAuWQb2KA8dn1fGaelywUM2i9gfrRPx0Ol1SuVTUnIHVO8NZ2xNB/S3EPDfuRs94d
LUEBl9qaAbswEqa34WsLc2XE2CX//7Bp1Y1IuiXfzkq0/Cxl6KoYJUYCXlfWoCYDBNUw53toCXZ/
lT5Gd0ZNCPpTlHWkQyy/YfLjqfvaDwBrc6cLmxmg87STDZiKe53ch7T2kiEWqBlmBMiQrf7U7JMD
qfVQVknCfGyAivKA8Gb/ilHAVuM9HVg4NwJzc/sIJ9Nd7yvyEM8/0oV9mveRPmqT2FiVYzUfJdN3
7NSI1pKf/WVvJdwUnFNuQlFuCYGGIdTyoEPzV5TcwNWyzYfsfw4qNBFITcjzfYx63x+fiCW1q21t
pDjqWPanmuAUT0sqiuJ6rD8OadK26Ke2nRo3ib73lgvDaAyQeJJhg1oGGluNcly6/BnOEp5GuNrB
/UjeFu6uttCvyqsIJWZMzjejT2Kd6qZ8wynhSCdROrN+hEAza0H7glWxICfSD/4OCsULixGt7nM3
lu45COrcYxkNzdOtOniLRD+JNVEJViP9jgKrSTqbFYCacqR4Ptq5NRiodXwNvNxeQQBbeX40o9ZS
XTzgkuh+jABF09sTDwwv+CHihvbTvbMUyqBmMXXjYdErZ0SwBZd9kPX+41xw74CiFLUlKDnJJJtF
+vCarue5gpasB04YsNVVqYeLZU1i8iY5iManz3kX1z4sFnZdNlJeRBYShUrC4XMHPTtS7R3eULor
4BUlKN3CdV+uJkSx5mVE3t3TNJW7YgfmN/qYwftbAVM3gt+byJxwNn2PB4Q02X1hkK0ncmhUllQu
hU51SKGwiJdaOheoVIx7aeaqb1RxuysmbYW93m+GuqhCQDrxFW9Rx5kN11IQX8aH42lj2uImrAJO
q0IB62NFhO0+3Gfv2W2SAs9ELCAVQRdWKeMKW/lUyw+O1ATJeR9Ti4IEph7ASRqSqjSnM3RKrG60
PYkvy3kH5uORTDa732s6vsHb+cdRzeotcGfCeE0C7+lohj+AWsBTQPjRWXBB1+ujGBa2J71zJzPm
ESckCyd3+8L1yFPqWZNOCEqWV/ljQirT6xmN8GBC9bemRcXAq8AV93f7KRVid0gfX+d7mjSPH+zT
qGpzKzd3osbBjjHdxs/P9RBaGyXZotIGkLwrz7QJxcym5eLkVaV2VqvKCWkYIWPs+rZm2sf4l5lf
BrlhWHwKOwqhQrtH0W12D2sdl/9at8VOJ3epX9i0A0hHq66TgHR8rS2vydd+0feiZt1Od1MDw7aq
WHFXEjlk6WV8k7acatrlaWsVFZZ3OfVyUYnvVj2fspwaLF4uWnpoTYwkgXesNr0E10mPWpcfGogK
YrrDMwWmFguRIsyOkMaa4rOL3HtWqA0hYvV+x/qK28zgSdTmBqD3SM9Ea4KGE9lABGjaP+1Y4MfK
nDP+L2F+w4lHW9W7qRTKdJFuxo0zknBeIh41eiFaTv0jajW97mioTU8VlXOCjpWbJFQ/IkGFwpoK
ReOCvX+KFr/qHuIpqvJvtaqkVyK5sRBueQzkhYYjrzCcwXndaAjqfMMARTXHaNUYmPnb8s6/jmCu
Wf4fhZ1cxIIHgywxCu7jnYEjQed/v2K3o6LjuvvMHtdysRM7jgaCfC6qu9/swH5AQ9M2hMPB7gF+
i9TY1YyVBg8cxY17A6uspBfZudiqPvVixnn7CPagU0xZ+6nG/e5IhPbLl0Kzdxgeoy/Tl08Ey+/d
uYUjWp9oSvWFwA5WdXvVRc7K/XB7nt3dqbPObhT2TdoN4avlF3W/jU91y7W4KDlLs74wXI5RdVvg
jAFvNOcIotVq/urnJ4BVOBJkVRIDdjPsWJ8ZiQwH3S+Pi8aVAHmhD00tbfCebGhlcDX26JqBNlhu
wwEmP8XaJF5imtaL0ApRVE8cv+UguDF+CW9XP4Eob2fJZtYcEXKl/MpiGH4B6yFx/Ds5ojhr8jY4
5zIRwSzc1jlYcjK8cQhLaUaxsJcTnqIpXsiioAvFFxLr8Kby/81Byti8OZMfKawwFwNWOEUHoTeD
nuN2KWZV8a2r3TCrtS8xQEfiTafGAeqvCR6lNoZzb+zJ8ud+AvlPC0KV8iF+0IuEwfVjTSfLY+9B
e+VLZCesCJyNEZp78BFcyYJjHyYSwwj81bjIXL0ZQrJkRC6TrgDUTxUPUSSW5wH3J+nKDv6BSXw7
6qjZhIvxN2aXT6oS/pSgFgCrKFbAYtXiXwodlXKs5MDtF0JqXuhOcE6A9tj+MYGYEI1Ui6VnuV3l
QxXTVVCt7wKc97IsGvlVyO9+HU7v0JRHEF4YURhog4vRD+XPOy2RQkwpRJETIFfOwHUa1Ec/CEEZ
qjxVgwxzCUUvVbMGx3uc9fX416Skp8P/0GtFlnpofo+Z97ewTnfJeG/oyksKOXeWI2FmHzfbUT/w
7Hc6TZF7yVR3ZMf1RsSJW1Pz/kURYaOAIWU4iRiw6sOQKQy/F4i5QwGWq+ATn5Xo3uuoIWX3uwvB
2uNJqc++IuTgccI/TIa6KsHR88NQhbfpOnCEN3aCMZtIKVyX/Lap1ZAu4sn+bI+w0lFfJTCkjNLt
tFBxxLIprRCufSOtX16yzzLemnQsLMh1qLVO1F7kTjkh3gf5hYyw7DCC2bHStYfG2gmgojphn5sJ
yL+EoDePdrWQmVd/nvsa+CQpe/uZVHaGAp2b+FGF5O0ME2dzTbug8CYWYJXmH4XpbTxBh3fgeKkw
a8KUjOIbkb0VkFPfv4Myu9DdEIIHYel6tc8a7emQ7doTtiBwXENzzhhXOcwEdwXdRjETHC5Q32aI
ozR2pb16PcL9YBnIQC83qjtINS2uyS4XXozd0h0nxJM7ae413aw3pDqTIU4XhCuHjPtgPI6tdYEe
fIAFP8dbZhAe5JatuCQaq3rqPSveJWMi+/T6/QrtT7g9XCmVGCSQnoFIAg84PbK4jUTgOjL6Jx5c
Sb9qQr0+1vWfo9T1cFMuEvD8B/oIbexAiTsU4n9HVf6MXcoH3wudZqnMSWQyJC7MmDQk2jD81VzT
/fKyHnVmDyiW/Dh9evJB6fOjbX71toST2FJNtxuqtLG5OXGbB5pXIIhEIwXTEQUyZ25NO4KMdfwE
48LrLbH57yPfIMVFAHTRDD3SoaMuae6hEokfOQqtd841UQm/l4BaDxJo5gF9bO4LtBZxnR7k7SSl
vGokme9XYU4a38Y+in84xKKc2cCy0+1qZ/33tZESPVut7oP68N0dg5YetXMyGfU0NTSB7FysQNcC
bm38ySKiWfcHLiKmxsHldbs49jpYX5ZQ7sX96mdqB0Bu0gyHqUwtdmU3l/09LfN7IQDyVc8YC+Th
pB2PWarBHBboJaX08HbT9SFvNYKveOMe5/RSkgcWa3UkI97GMWFjuaQfIPHKTpEJFlhXJsz1CZGQ
fOk8IptRPF0UTYO9yQ4WsigY2LdUiKbOtQQfjIDs60kfePO2JtVrYZqmVKRUVxircv6jE4hKfYw8
ffrTw0E2ll79eAibXQTTZgxIs2Eky0DexMRz8sNXn3TaTcquvpbU1aX5pNFBil8xA0JQxLePNv7v
IQj8GYpaCtCdpuzVSs7vwZjDXptxTUrWfu55FugBnyx/g5pqoBLs0mqjrD5WlsEAWi+2k3HskI82
T6VST3qGwbq/PazLlRe4PgKc501ufX4vlZ5hPLZh2SThfCCra1NXEU4IzQv/6Kd4tKqgawe07zHO
hION+xNqRC6Yd0mwJ+lf8HwnrAM0P5wtkBr3CidSz7pyq+H777PLqDQeKlz+Gu12E6/wQQn70/l1
JxNV2O+RBErlnSbvY9gTYyNHwbjsNT0dGDfyOofbcVKViMfRGZ2FxfDt1KtQm+ak4hW4CnLTpdQs
b+iOHeyr9WehtTa8+kM/jec6ANkrtoa+PTx2AH/YjFOpk3JMWiWsjCmbPs4a4MbqEVS7PWtGj5iy
X82lmcZ8QVmF3V7xIl4tvVktIixLBYeKw1cfpMRIiV8LeDFRdtKn205uvDNMMDpUtgk+Ik6pz3gt
v4VDRUaf9UrNYy0NtuBGL/v7+wONIVuUnx/v3O549N3rR8YwJLkXILFPj/egxMW7ohMG+c5jmCVo
6g+eQR+5xlNrMqg7X6i29feENrlgV9p+cjajLhb1dGFVYLHiQlmSiO/wOLG3ms8rjExs52ju05yE
fFKTveszUus2BcVRgIo7PLik5VeSt6bFUECj7Kk8d2OIN8gQxBONK1uBRzXeAtimeopNVt25vCQ0
KUWLcNmhcPzbz6Fc7BmIySozw65wyc1atuH6GhbuFBtU+cYKwMNz5XjMaVVW3xmesyOPThpXKkJh
op13zMptUjFDE0qL+1KJD6D9bAXCvIiP9AaAodoRTb+MuoYlpwvokUdHeIzy17AxS2P2JRes+5mo
40w/r5OOSU52nw3A8ZajmwBt4cUVGb4yvYvLi8u8ZcAt5mjUGHrIlIlTYdiLrxplwPrObjfucsko
5QImbh4aAHuE/HWIYp8s2CuAsNsD4uOGdAxRqJERVD650NcS4JKWQ0MET52FcwM35lyW0FBdNfQ6
H1uSv15ifOyOlnGugVVPx6jKf99NduASLPytzvjz5sZN49KywHjlOjyev9amxrhtRBmDO3Yek9uP
qPv+hF3cTUeuQD7SoHEHbCBxBNz+y32ZbRDbXzJAne4HC7RsrcLe9Md3II2QMJo/jxG4a7WJHLi2
OoaWm5LjgiYiZVpPS+HBg4NRgM1JG02Luy0U9HWVt7a1S+YOwz8roSoLwKVzPbSFZiqdu1OIY7Rp
Yy/oh7QE9KLEPyqNaG+5/+oIeAFJhhYffdPyPk6HNhghQYhVFCn3Md+Cr/ILeWVxEv3A9aaoB5DK
LszysB3xAcInn4X39hTTdOySGOgyqDTiqW5/8rFJBcm5KmO4Y6iKPMBS4P8+K0s8icJjWjB0MrW/
AdUghcBHLNGlqShg3Qd2TFV/cittgqRX6ROEvgCchEgoxZ9UECWqxrWzOqmC7w5MmgriRo6YmFiL
w77wJNlcoGEMcVyiVMCuFPdMyhgajp1C5nR0dQzFGIl0dcWmwtr317TjZDA8hNXPQfK0g/z+OVo8
3Lj+/PqkKeyCUl6kV2octSWuy1ypVt9nxUeYTqVIgjN8E3uMm3tqb6RR7odq3hITqJ1DfIOxHCSq
H169ioexM+IneFnvet9L0knsFhlY7fZ3yB01sRjxZdElewLZdiTkUCkX4Uk8Aw4W8HaOmX6pIfK7
3vu/pmWt9rWMLj2qkoQBttKvUgaKleEc+GJGOCvD36XhIy7imcwhhET4W0/HHWaAJdKj+NWSTp6B
66086aikEl1SHxF98yQcJ1Hx6gItL7LKxke5vEiL7NcRm+dbCzBRBA6vzg5Tq+gpqyz3pUv/JCjh
t0bn+2S1gINl90gixix9lAdS6kqvbIGkKw86qqf1/rw2nQGL9+WOl12F3lEptkEBN4cmA6DiUBgX
IDAHiVWYsibLKPImwu2MRTWpt/qQ19BTEmNP7DXEaLP3nCqjI9srLbaPsKp4CCcVO35SWl+yZoxu
p75L8i2PDW5aGwzVSwjBO6N7lrTEQ9C2z7m5SUKGqbKut4qPJ16AHH0uk4esPxfl20dEP9DxnfA7
Ro1+Wo1mlX2DGOlPb2kcK1Whb/aC76FHzk/DSt2VW7l+vNE5MqGUrdw1iVjb1WEGW2mWIBw3/QXN
ae/HtM5WtFk0pXwXVP+er79vfiH2PJqcnNkTN3UjCpYf/qH/Az/kRsqjFnozVx1nhktxL/N90BPb
VhnpHd7hKvdN2D+dKopnITI3NgCwkGbjOXyKmoNYrXpmI6+v28RtEwx7jmILF1l8/2DT9zip5tUU
yVzj5TVMdyTF+TRto463977puPLaHi6fUv+wRBB1KgyhXCqO7u1PgPLuhOD7FVUCZwpjLIeqYwVV
61JPf/MsY6L66cW/kssptS3S4QbItNdb6in+/CFIM7spVcMIUkE/eQGnFMxULrr17cRWF2gV1VEm
5eNSScbLm1hJUtzg+RyttPXU3kWzgXh5fcHXJU3svmu62RmViqp7SmU/r2/wiUKjW3jjvvvUMdEY
qJqs8LFrsPvWCISftOjTw1hbJVwBg4JC5+GZvksdle7ey1vzqpkTOuhLF4zEwamGDQCcM461HShD
cLUrzLvTbAZkMrNLT6yzLxXtDuX24XaVyCYXl29YbBIILThyGEeuHh0r+SESIu+4gwal5ew1syk1
gndepd0HXrR57XqmjzIhSTnij0YcwYVIU/b599GA3yJJhm6GetIMB/tUmB+xMfPGvvQqKzXU1OM+
ZUfEr9rKo5mK4hNMiHSqi7ryc8A9GGyxkTW8HIBy+3TI2Bpr1DMuCp1FQ9xoBrN/i0sZQ9UuAeTP
4bTWDXq7sVlI9VaO3UinOs4uCHSy2av5DLk6e9480/POcI92GnjmW13xc7bv2Z8uKXroct1JQqfU
IkJPlCwi5G8GTUCsm0kZXlotg9b7OATIkhw1XAtLyLxL/5W1Eosoq1r24xuPE7FXYcVc3SpDrx+E
dY00z7W5MrciA6PpOz+KhnJ1FV8Pkv8dKP4jS0hFgVyEOVSHMCbH6Gm4rVl+A38vBuPCCfD7+5Eh
pHsxTIHLDzDofy51CgKm0jKmNiYOlD3C9fkCO6B1+bixq48Xfm52pxLYRGou0PcbQwBguzK37AE6
QR7a3y6TiLNBNeJwZ7wVzOKzKbXoYBIAP9wnWoMqqj7gzXD2O1DVSzqU9c+W8gJYybMxFm4xPxSQ
+CCRiQVCJELDZlrpWDj3hLhTNRye37QaXkTL3spni1d21fK/t+7Y2AQu/EE6YtlE/bWoi7bIGxQX
LqRvITtqd1g4IX8KZ/zFW+m69yWzFiV7np/S83BJdwD9AfX5/5xEmjgwePdWmrG1qS3RYoDGU+dM
0EvEdJ9JPItH/KTB9X4TpxHda8P/5r0yNERdYbuAfTfe3Q8rJGevCJxHVkIAA78oGQzu37wFwbZE
6h432IGfxfPD8jVA0ENRejNIe5caXQN/QKXCdgPiwDgqZFZeIlxslrFcUGzfkedGf3x9Skx4fd4P
QJcs/O98/0w9Jgjhmh47ePNa6u1OqGLo5glM5vkYDIbKjZoKv/QVHuSCpZK/ONpXZN9qLJzC6MHC
8sU0iHMRu/SP2ylVcVRB7Ne7/FG+InlXbjaa/CdU+hp5W1lhU1xku2t9jbPMCc/WAaFWnKuwzXlS
1+8pSsbWljcrwTOmZ1lknBcthsFAde7TULFuclLHWerQdR3XZR75/QTRbAWy3gDS6Zo8TxPLELTE
j+ZAoRSk/15mFWStK5N+Yk3/Z0LNDaeATsUMIhRpP8mVGzJV+Cv6js29kaX9ded2iSWLIplahEYP
mPwVwffkIXkCx9eH82srf095+fWiPhzpermuh+Evc7PHnJKjw7BPoRVD9V21D6O7ZJ03A0slapaA
1QhS2M23Jr5DqIO5mzjQyXAPc7QXV56yeTR+K2bsRcGfVJYr7QUY9FOI1XBuLlRkPyuQPvehS+GI
I/es7iD7jhxselP2JnKENtyYx5m4WusUUHEDFbmHg8C2zzP/QcoV8dSR10nZEKPv0M47p4+JCYF0
F53QwBvLO3I3hDjeUtejpJHdgC4h3sH83YXW9pS632GhVeIKYLc+hg81EdrR2ArW8lIQx7FTuhti
zp77Gvzw9fyyhypMZS1umwNjbjS57MCVXI1nODm4mFuZzLtLDovVISln9YKsfvrOxyA24jh7vLMk
W/W/7Cl128wh48M+qqx1lbYwRu2Hk1+vt2EqsHejEjE7iLNQBAQIVWerghUhG/CzSBXbfsJI7fLq
NprOOCC/zIGchqj9J1mhuYzVN59BtnG3O4DSwoHk+QOHrx3EUl23FPCZPHroWAcRqVhKjtRZKGIn
z74t7n41qkCrPmO9eK9v1exIfZE2UrP/rFYuZieqhVpepAH6Dg0KCv8GQp1a2PPZfcuRuEDly3Rl
58UDrTTMY9sMGnN9I+33Bbxth3O7cJvD+NsIBJBmivNugD3+8GmkYK1kVwwrCWlB+75z/TfqQrWG
H834+Bdf13c5GtvExX7bMPIQ1M+jWLKyGr+ugY0lgdLdywABm/3mfZcxA94QBttkxlJKKih33g8m
pM8/MAzmoFh1g7MS20jN/1IRiCBQ7HuSc5NoRUQywx08Xjn0KWqlbyxW2BIDCW1II3dg6+vwGmT7
6v0lD2HL3mMBfJiSMUpOovjZ2tw5wnNc+rZVEIsrpZIcIHAz181r3F7gZSTDCL0DSHODsl4CN/yO
hr6VY26LUVNZoHMpL+JhZAYHU+gReud/72dmBNCV6lo1Fky6BlMs1iZBEZJbvqDnG+Rdl0IDMjDZ
eFALFb9cCh6vVXHgGFMzQiiTBbJ3anSwtFDzQXLmSpqzIYwYeo0p/kiCYWXVPX0fP8tJgotBl97h
AfBGVUMLKHBYN0uQ02OR+kGSlG+tc50tudEE472koOIudtNthy4QB+UM30cEg9Ar/72A++OyCeob
nWFB1lDPlRD1JbSWkNvDZdFtidPTg44EUFq787BLea2995hIDJHOFlc/vvX452BHYXdd2pXHKXU2
LKZ3/ArcKdh+koMqt+sPWJJjMhqkDJTGrVJ9ISUOZ2ou4wx2Z9KrH5mjkcuGgsTmVu3ZghtS+G5x
27bRVOnyD9/+L5C+/N7hpy17nUUz4trvgq83RTP39gAwswTyo1a+ime2tNmD/9Q1BtwaqmJhzeNe
s//MTn6cVYZ89M72guSgHkNLbkC6/59VVaxl+avR+CQk7rl8BrFJwDjSadQFqTMVPAXXosPF3j1b
RuPhagS3suLxc0+sHFag2yWteg/lysTRjW8dovOM9iyeKWDJErZuXOD/UUbHYlJsfWVWyQHImIuE
RWo3Kf5CtG1z6rPDnK6hBbrZIqzJJGnyr4WJWoA4pNehVF4+z42YHwzZQOG4ACwwUU+ipA34h4Cq
CPox6gVWCmXLncCfqC4tU2QmsLpCwIj2E28dFmuJIHtKLAYtdnrJZAKpaBgGzzLOGIE6UI6dZ8z/
b4i72+vwPIMy3lJYHrs9ak3FBr1NAYevOBquzmIIoA84zoD7gn9YwqGAgzWtTrbbrv2WRMFByWIS
5TSP0IvOi285zekSMFlJmguLlyfNJ+ALXEDfLC3yzdP8pB/4g4/okZug7epoDzWwifzpeEVDuy1o
Gu0+JjZgPOCZZPItJRmNLYjmgC853ENunsuoJAIUhpL0yNfM/6dmlLaK55n4Buk+22TYCgJw0IYb
7Fq6V7CF2bqc4mVD/AEiyBW1E6e5605FgN/7u+lJb4gAf47Dk+mosi83VzkCgfTWvi5RPi1Lr5fW
kbrHlHNIprdCFQEAvY9KZBU+NOY4nI368pOB6cylEJJcnCCakoBUliKsSOGBOJgYjFganFrwr3ZD
wgwUao1iasRoTBhGhwsT4m7HG3tprKdkpHN2+z0sDCPy87imO1jaSyPgELJLLapgLvTJG9yIgZI0
wiOhiruWl2MuqgVQ0YtgWky3DzZzfkHGxIMlYtac4/DE3NB0+qzed2/wSlsUIJMioSHXXQ9Xtvlm
TjaHdOT0wgcIeDzIVgrZ+J4UQSER1KtQebA9n/pUrwGanBELb/645koUg1Daw4oE9bL8OJe7nli5
pZa9JMlVige3SspU0SlP7wRQTB/Ak6Jomd14F4gF57rqGrUnQzKyEfEqW82qK+ZE0yeKMfeCdLK0
AW2J5hf27OkkX01aQ857WgK58D95W0R4NMWPtGg1gey8R8HUh33lVWW5hjxYD2o1YToBPp1YRPrm
jTv8j0VwBak4/ZgLX3UfFDVaoReHb53oN4QzVX5Bx5uXM732Oa6tnmhuTTWDq4bhYHZjp0M1HL7x
fyEbeVTqV2GjyaMro79xOLWu96F9JdqLRIZ2FwUsVqDuogl4yYxciOZjJj1D0be+d9QAA0vCLlUZ
uIMjCnfqh3nOkmBahx6QB3/riuV+6oN1jHlERZ79aa5K6gYKpST9l1tzl9Z9LC1Ev6SUhJ3uO4VH
RWNt6fPpW04RtKXmmhxZvoFLEMOKqSCaTz1fDk4HPa2jXPU7fiqwB62q7Gowv9i/QcFVQfkh5iOX
fOaHlLC9Fu3OpG/s8uFq56nDY1p3IVD2veLu1egUIboCV3s1JpK5FK7chmKdTBHB0DVQmg3nLOvy
oSbh24f1kddgzC+3+mHlEsb4o67FZzXlq+PCYLp9jjG8K7s1y09zzgYm5U07KC+DblBjpUN4agWY
+CQx/RoMbhIx+4UsjuV6Ujx1AkqsjItZ4MLsYnr5yJQdKwIW2Lo3nBh+Cx8Be8+X0cTy5shaaPz/
DLddzKMdVx+6ats6iDSM0kuFPu480jxkyDPW6k4f0GjBy/41bIA+Llht5VQaVVncafUYVUoRsNtB
FRavisD8JXFAvIx+gHdkvLOos3TgVGgyN1D8HmSpKkA8lgAQkCI2Ixrg7afBYzgVgs+7e/iRFkqk
klZ4LSPSpDQ0rmx2so5C2Q9BjBQhhXHKG3hta+svVxbkzq9IFRvqpwIdeUqih2Ha/btpZAOucu4o
z0Uqh30vTEqT8Ftz8XmQYmk/4T711swTYiHpXIUUUJb+Nbe3D1Ft0C4jPRbkX4C1RJR5be+lqkO1
HPrOWWHyWNWwkJ+zKEBnRRVD6dxVaFI8sfqUMmxGadA1MZg2dTcNp/x1CE8Kc++2lvm2Bg2qEYGo
K9vnyzU8U3298G7zJqOyZBaeByJ47bp+MUzjWuVMxhyTsitq7u4c8abf+q1o+w/Tw1aCayYEltz1
s0AtC31h1RdwD5LdhMeXhzzfegqhA+vRMQGOufL+763TxM07pKqMoqhQNhuzkFekdr8gSy6dWomQ
6+u8WMT65SHN7BCHYWJXW5hqe411k8e+NpLU2tYRzDXRcu4+d9BZTeT0sDLbeNjksvnvZYzGWrxx
6Itgjcx3cwirEW8ybODy7lOu54pk4EqaKJuDIy4sVIwVqD00latCygtWyuiqxwxIUEuSm6iEV1kj
Wu4X7TV2rUJSlsYlL4nl/mFbTDq/kTlGr+7DOyZlAXrJA5kqmzY8zCw68xokxUTU+mpblAg/7aW8
uYEDeWAQMnj6qwQTnl8TkbV+SG1LtHYQlBWBzh4zrlS0xRNEcE+3tD07mXb3ncOdp5ZpjbKpbZar
FQyFUA4bGvHWmvDEiHRRSVyer049JtovaAt1zpp/VUe8/NUrxMfTje9spOrle36KgpxA8ykvrWxX
yWRr3DXfWuCXX/oLzRG7Wc3uRXOswYtPn56RvjdpElaMwLIqzpcrIBM1nvbrw0sze6GfsJ9B+l7Z
7y7iIgPF/5YI0ONf8T3NO7qplD9Q0g3l1ZbG4SOlx5UcJN0N/jPS1za/gYgwhlt/g0gyQSEvMtFt
XCVzPMWeJRkW+zLkbpwC1jmymhNKeSjYpLpOaWskOHTQsxIztExcBzYOsMV6R3zaoQgalIIaqOvF
PXCt4uaELc01XwyUcqnctMzWe75pzyIPobqwr6vHUO5/TWuXl8QaMvlGcu9d5C/aEqq5G5FE0cfC
hVQ+3MGt++m36uoFOuv99QffcLjF5mggsBM0ntaRdqT4YJG4uYZS1T7O+HUHIzKRMvF4762U8ep9
yOEr/1Zz7qdFILJZjRtIbJc4MvMEoWa67PK0dPt/BiH8NdW7zXfsU6BIsUZLA5nQ9hXE0Fu3T7zR
Kz5UfM3GzMF3XrbssH1HIcOqnm4bHlSQ2naZxFwb1XlN1eHf9CIPDuRqvbwWpJcEWznLP1W6ZCGG
7kuAxiObSXbES9j3kpQ/YYxBA1cBCYyI2A5IRr+M9h7hlcRmb/24bEy+YQSELGNooVzEA3Eg19fh
U1eYxyCRiqvWqKqtDrSSDS/IVf0fUntORNO30DX0d0r/Ybt3qCqAmCiBvo5xqVFAXxXNSGr/awQS
ZcyLe4njgGv0HHk3aYhRwH9zJefq7HVLfH23mEtjFnv3yE3/dA5uRwHdWjR2gwOUtgnoa7oYWmH2
cvy6/xDQU47rDD0fZbvD4L+XgvU67WQLvN9QRawi308Eof8K9IHnapDczGy7yyFPZcNiCPj5C61t
9G9tYKZE3nddK/QLpl8XBD72wuxfpOOc3qhjyfSS8NjhNDCn7eJynUhvfkjvQApMpTRxqKgjk/Dt
3izWV11cl75QCXqO296fRfM3fG2Q7Fm8IP6c4mxasbG8TmxosJJI32a4d4J9TS9Cpw8jlCS5heiJ
p5wyeWfalIZz8pXqNXoLf7i9l+kMYcXEDoLLHlJBdPFspPWbcMooVwaeXbwk+/rxPkxQSQLIEBGR
nmfScNhO57bXuL1V0BmU0Z1igufrr+NI6Thh7W+n7Qm+HU0LYgtfvD+s+ffmTM+IpqQuF+9RvfH6
AY/TSWedNxJCyxNs23SPfwvPm28VXqB7igOeekzDkQMHSwuWNMAuN8PK3ERr8mpXqD+EDsxvyUXB
9NhjVfVfCop+tPEH1euZJU5GgWCaYziGra4+zGu1R7OsZJRF56ZMSS4LxyrrR4tI0kWxbEYKg4fd
pU36RiasHATwa829NIlN0yw2ajuTHITt9YBNs7RKEcPw2v/a1gxILJ6GHJsgT+q7hnKzxY80HPyv
+oHFi1P+EW9RWuGoTkmBFi7lowKSI37y59Cl6REzCvEZkkfBwUyPYXOklhGBsuExHYwZgSdPdqp4
1g4H8Y5dcgEr76X2no7QgxHQUqvCUWQDX9f7Uri1Jv2SnCad4YM7hgSrC3jq7CCrMSB0Gd+jnyOT
1bwR7OQZJoL6HH5o7DKgc6n9kEqkHXW/tL3YkxYOSO0BZaoLezHQgcNuUbd+m7nhryhxEtqyhRSk
L/WFtOlkMkmJtVfi/2+dBAQLzD04ojW21m3MOnUXGCq5Cres+KfiKQkxwKwkpq1iOcbr3EK+p5VN
nU7LqsXNbpVE/lUGAUl4tmrqS28sJKn/tsGrcOzy77wLb5ZvTUmJZkrDmVUaBUXV+wsU+nXJ42pd
/0XHWRTWi3gKr1u5/R19JafCIqeJlZGEG0z6bhHxxb3P8gWINsHI0hWNIt0Tj8hv2zMefNEnPmfB
PDTO2tidxvZA8RV/0gz2rs2W+fGwauSeFNFOS6Azi1Ysh1/P5FhFhG15oewrbB+YIsEkQnIe415V
Ci/e/tg3RhR7nI8E3o9ozWopSCRA0xXgwISj2P5AMlW7YG6sDcoAw744JOjKtRUE6Q+jpsD8wjCH
38lSjOuoXL1sXHgdJuUThGaHfmWU/KZJX1aEhyUH0zoeud++yBoLkjCelfiDFA8oWyv7ClnzHNgR
rTQzrNp7ViNqpMS/mh82q+WEMAlXRQ0Q+rfs/l1sQIYacYLDoziSwKOrAwmZBzbppqGBDlCJ0OzE
lzZxBmOzQHPr9temD9rXh/nzV0U+et0vhoqr9p9BV6DbuHkKDWO2BG6Bsl59TZ0bYniuYD8HkrQ0
jOt15dMGqZU0b+BcVI2DuNZKuxbUJmFqyo2z0HiBgOvv8s7xA/QBSmgnyOHncZFbeHC8ABLUgez3
7uXcjg0henO2itrbPUz/9sBa0gUV7e4Zay+JgURkpwDXEkVJuwT4Mor7VlYCZQPmE1AFn6ATBLah
IpwTA14dg5m6LTrGfl2ThZoRJQLpIQbryzEcVHziZj6uCnvlIkDF9kBMPc7b7c7O6IOVwhQARp3e
yM/0XbD9tRWLV9eBMd9NidGKdt2JT7dk/l0zBcfCUbLOTa8TzLVyQeDWKX+QFBDK/zLa6yZBLv9h
bz18sYDtxDE0PurCcp7BEWdI9JFkEdbVEw8rjTz0vBs6vUpUwtDJiKTSSC5P5S0rfgnfapi+7ASZ
zmmwfDIrJ+vmKEvLe4+ULaFbPuEcZ3K4eCf1qjFmq9TCwBhRRn3VttPK2sJIf9e/w2/AI3lzUpZj
nxY01mX13TX/2r5GncBQYc3UvyHhlsSS+kXVKXxc8GCUaQRcdLBakUxWCBQMjUYQeiBD9Ct5Qvk1
jtIfu6QVCfcwg37euRenOAGqMvLu0WFbmVMx5BCp1SCROoYh1im6zeb2c57eWwVGc+KO3EEiBGDi
ivfCt34Q5V8zHZZqUBWYMbyYcLf4TGiEcSEpCqTWtCH5S3AWFc5/9laquShIahE5Helsk8L6j7hb
UOGFbantsYw8dnpRopMwVcP/B8s44orC0BzwEAnnqPsuCTmoVP8sSASpA/DxfJNmAbOfRZH/2BzK
JZgYDn85nJFGfs2ZnGIHx4bAwMD56aL9CL+kdBrZsrp6DtBuG77Ha/1SloK3QTARXpkNS0VuBW6G
prosMrxplOFWkEbhajujkQHJIDQVwCrFiWh7khFHeVAaitbHSolSssHLQxGCTCw9jJdhRiKI00kR
TlaigDNGCQHCfbqf8TRi2CwKjkGgvMabMprSYazW6L8mbu1Dih31IEk2b/Fijp0=
`protect end_protected
