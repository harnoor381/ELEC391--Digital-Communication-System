-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
mdQUMiXC4J71B2FOYW4uEXAJE7ta4hg6tn1rbffnRVm13iyiYw75jrFWRr+fToRt5Tk3O1MHb8Sy
JjIyB3hjA8pCekjiDfvyBHQn5beDEj/z5uzd+pm1G2ThsQX3B7QD4Njpcy7xyns1Zb+JU4avG2Ss
Z/vFhubdTIEEMGnVGtlIOKK3nlox20w2rEe3jHZAEo7b10c7FyBo8mmIiM3ekH1WG3X1YpgSOEbJ
YWK+wbRXm5wIGksbbLjTiA9+r/pI5hxdUDQOBrgnNFJxVaLtm+7wXpAWU+NF1oN/H9XdZbr1cmti
AWyR/UuOU0TWi+Idbtu0bF9N/Yym3nStjDC37g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 22480)
`protect data_block
2v27L2AfM4k/K8CvyJ3JNUjXOOoK3Zcedoq8FVfVLUsvar0rILT85V+FKSkhEpxS9X1OyUgi28fa
BZdCwWgwjisONVRFUnEJCZqxD0XGAJj8AhASTTX9Hclko2Q3ytUaJi9B67PwWQKvC4omJhH99TUf
ZUEURjeP9hnii31G0yWvV/7vud2yvg+EUQedKBMe8ZR/m3XELBZL/GvVV2Gbz7Cm+/GZvdsGYFkL
w4POe5p6pna8jnPV8lw1F7PTmebNZ7L9b8n/VRAfYMbhOWDjQTZABx1A4iu/gvGTl31ix77u/Fzn
4NWOyOLZt+oJPDXfsLwT3op+T0y1VCQ6ZEk3iKvdq8o9cB6yIK03QOqGCfgeMxQ9Pqw6bIeFajyk
CCxQxPZkZAFURil5rcq3M75W7KNryICdxCyIbfI+ufHUv5iSFSz9iKUXqHW6KbwwZFa1ZjTqe9aa
OQhZkEN2i/R824liEFXOfIYELalNUeN9Mdn8R8Uzr3eJtQE4CVNeXiMehogDn43sKMArTyBDRNcg
W12C9QkX+O0zHJCsHxaZxiGlUB11sckeSs6LQThpcBPcSmgpKoUOOgbzo6aJc5LBcWRwKLjKajKE
ha8F/r4XqWcWpKmmovBkhfbtSAtAoJn3qQUwM8pwayYVNpD1FghXvTarXYItJ2tjsuWEoaMvaOJt
XWzMi1GVFbjjfMzh1PC0i6rE5Q8qf01cq0bT0dJ9gsA8ZEod0ju5JVeoMT9qsFNh3dv3O4QMLqTo
ZpejWQzPuv4rKsxYDAUgFO4a1uF48cGP5nznFWF4ud7XBmshpYH4gAPf92R2zc8TMlXFM7HuzDxI
oV95bWt5TNHL03X/WaWahunxv8AItZFAgPk+vdEzcdIF+XIbv5fR51x+/J52JQYsgo5+C3QWTWMw
N3rtCmMFonJso2Wp5eyTL/CDKJQOp3gr2FbDiAcb46DYKNExaudYtoyJZRGO2OPQALRtjNApzNW0
VXeitRjVf15/V4F7jmMmOjvr8AAVS4iqkHpBBLd/fJ12dapJnvIAqroVDyencuENQpqHXVFitc1e
IJZBwh5pL5VmtS2twNswfnLtBRwfGf11QMcF7ZJY8DnDEiZSkmdiXFQrhA52EYF4Ep3oAZ+39kKO
d2R+fLC+6Npq7p1aXkpVKRIng6Cw4tZ5E9SJO178/qKT68ZR7wBnsU5Sc80Jf4HuxMHEhlFMwhkj
fFFCQBOuyZwDnOi+c5rH9pLndN6lc2PUyNwvirc6uQiS3SRZ0OcwGuyuj9k66GgOzacrrFZbY/7i
UkOAF2WyFeXax4leWeiQB2rHf52kowyncM456UaEf1cD6RlrZ2PRj/7O26GKjGPcssgWCoowgg/l
hVHgErRbnzUuwqh+sbmnNtMbl89R/Da13OCVDwjOdFeacfKIBjQuBF1ECOoTg5FsxXR3EFFCD7bm
f1fGNT6W6X9Q2Rkb9HRMWUZK0vK1lqUKV+QUMUJXr4wQxU7DP/kFScJwEmNXxpXy4pohKCRXlwYu
sDoGlnMYAnCUW9G1tj+28e+ygH+s4UOi/7c+sNgWRRDFPbbA5ZCzIJIge5GcS1CB1sq9buLMn73M
HlKQ7E/X8rd4fPwU2h1fhm7dRwleJzlKWzhSqZDKYI/rbDMKIznBHkaa09aNBrnNsYPKAQz3FD0K
L/fYiha1a5GrS69FKcoY2o3xXrJHhlHCFn5rz0zvSJ5lBisHohMLgJLr0avnRIjnXQAIXbUz/73o
mWOqnIDsWQBV7cIK8HxxwQUy3opIquYTjvqi7c8+wW6BM5suYje9HVGZv759s+phmAkqOlKwou8i
c7uEFklL0CMjXvSiDo63ZEFkIYSd0MbhjyMEzxrJ/ZC+EWjlCVdjpBbjbN4y4W7KsD2bn63ioghH
ft0e//X1xeuXMLhWHlqjLOTc/M2cOOVfn/6CTuOUr1f3NdXqOU51yGamwUVt8prp0F7eS2Y1wKr4
iB3qT+gk4TSf5aNQycz6I7pTYMxd3YDcsRfw9cIxpuecDVxULPW3PX1mO8Cu9zi+iVZlRIW8bOAl
WkD4BP09rNsjGnurgoO7LQ6jiTSIr7uKSgJLSks7De9lfogXJ4Eja94MtD24yPS5hOMi7HIJAJBI
M7P3Mqa3ImAn8UZ28TAcDd7azbZBdURBfUtz7KLDgocrKCiPdUBnQZ61M8LBz5ejVCyTtO+pC35f
uwBhf54ImbX6NOj+aQDT88+yLTclm3WqplIk7E1ZuUkn2F45DRiUcYoVoYAJuZRHn5K2aqdCC/67
AXsq9zs7Q8/tTQkv7wUdR2NvQpHiTsbG9+S1nPEIBsbtpArrTk9zLuRn9lNjxYuZuJ7c+IBQSsKt
BQm0T1NzkT2QEFvoYLUBG9htzqt/8J8BhJN5Z/9j0uPd+bpTe7lGL7PVJXJPdA3mhS5uNPeLm7hS
Zw4No7goFz/FsrAK6oYBYlslv3PHyTMwG4R0WB6dfL4KWwIKQaxCN+87ni9MU62w4ZzNE5EkmiNU
HycrWNEnlxqFR1Y1D/x2WkbCjMFL4B78RbY/Z3XLSOl8ygxJSkLcqlCAMfnFHLXk4eg1r7Tkzboy
X+BmvI2ArF9O+XyuicxZY83O4duIh1DKVi6PUBy3oIs2C7Bm0VJVccyC8olGaJgcRHvK5Nl+Itrg
XlSgiloUhmcUPbqDO/MyW+kKv7o62Iu3yWtISzljXE2g+62yg2jL+f1wLbw98T/361xXbL7T4O0v
q/uabMgWfVNP1J2xCJyuKXFvcizL6P/5mV3TA5JBA+wuNEwINyeD8vdegdfe+4OTRj3pd1zysrRT
5U7MsMc1pvIEQYV1I+2VfihqGfXl9JhptNXTygCmeg18Alsyq6txxx4ldI8CoW5JawG3ngixE0Vk
Z7ObUFFxeJAUkx6jJkh8t8HPTjEhKkKCkI6nYUaiDvO9wv34wb1rSzfHLpKnwmBeQZDsPmI+c1GD
nEXFTd2ROv4DK/LRoRVkOcxMqRJlmzO5U2B5vNlei+zZYNVQ/nibYsUY060FfqB2JI8w781XwP0b
KRgD2Cautjtd6uzBSk74PheWeUqH9Vf3mk7ThZ49gUxAwHxYSviUGABn+YsBgWfZpYws8sS24v25
K7OxoUYKYtKmRBINfO+DHVYcBQ7Jrn/GSl8690KAswDam1m1b07hhIUKrlctdP6b3z5IOa0TblIZ
OAGPCCAfavPpri5KG+NQKZ27qJVi1E/XtGL9IZNA9BXAxyGPHvcFLCcCagnvm2VMgnazY+cLVxyh
xhh77sKJ+TgVL48aNH5dHNIoFIoTEB8KDA5xbImPvjaI47l+sqTd26pA2UPkUx8r9dzNPqD42IG0
5OMWejg2vkM3mraNsrWaU+IKYLM3tdo8I1RLOrO70ojt6BcWvmZRZH45mQFvbGvazsIcEzuAglvF
0E5iOab4xsNvbd+tnnPoQJX6DEneUJtAO0DJgUBUl88XkskTl26J/8vHdhExhkHIvLb48R3DaE1k
CqkMizC5K3hQk0O8SgUEloY+at28wZyUrZ+dh1ikNK1Nv2mePXUhEeG9QWzB7BIJ69+UUKOrm183
NqcFo52TloSKLlPV6NEVeBNKugR69HkeKMsEdxtGNQt9f18v7BOCXcUJhja/7OKFbZFEsuYtCI5Y
A3SInM4vrOM1AXRfGQcJynM7MpFDtIZzdd90XBl7LGhjQaR7J7U3Q+hv8FD/ufcTIXwLSLWFBg8U
jVRb/RMnHLGjJ/F/ur/i6KmsvOchjMYJ4YO+RxKV65qUN13cW8uyRcRvS26zOhbqiSgvffbOF6Ii
aqhQY5dtiDWtklGL1N39gpcRIdKMqgVST9Of4k8tbrEMcQsOKw8hrpig+ImpX3oN8eFGzbVayelw
aw1EKeX5urtISZqJThJs08Mdf/olEHTDW0UGP+Ckdq/x8mZkThrBCETyALYBe9iBb21iHmUl3BCf
NymxVEPsFiAQmB5JCGiM6eZ0H0N/s6p0tN52KBXkrZyf9lcEgMH4QLUruRr45t7sr3arhUNLefqZ
tKfL/fBwG7TBbwZptgaEPwmAYq3nv4CQZWtxte305Kn32Ndm5LxEeZKycP41R6G7VpNj2t1RWDE/
kE0cBBA8N8bxmeC8i167V88BmyabP3/ikA+PtgM2SAbusnzPT1/BfS+PrQgNg/GbHpSdLoqwOO+b
eK6oB1SUwUg9+KzaZ1lXrchqMxgBmS7LYJHTI74dwXu2qtEw1F1PH454C84uebn46htV1oK9+nKt
wlNvO+t+7/vOptSOaVnyFYSvtDCz7yNQVssZdWM40NOHeeUmtnCZgHF16w+u4T+Htsb1YR1/pDKw
75OTlpJfVvhr2tt7x0Psh15WYelD/k3gN2nlGk9EyNxOPNx97qrU5sYBjjjYuKtB4FCFrYAnQzdF
W8x/zsmvGlJmi79zBpcxW7m6zNXLeSnGFGTTLLHceABlErbPhx8XHsYpMUmmYjy7bEggZujSnl2O
vy5VuxytH0ukI/tqrmvuSgoZ8dlogtJCjQqJJfOKgfZDdrxRaH3uW4X7GPaCBxXOsMmJEn3jJts8
Knm0ziDT3ssrPLzn3kuOxqjv5kbXlL/t4lzF165+A9rWnRuZmUvGEjYaeH6KpIh1kmPEjEodTRBU
ay6lm7kdpYzbVPsHWb9owI/M3Cze5DkjCJRnS/Gm7OEHGDDCJ2EtYGSkmVdrV0k9VsQQGUh4DU/P
8XUWECdQi8gzDrUkJpD5t8Bo/LJYNwiWQDfSwmE34mM5nrAwWNCFOwW+rtY2IzqzPlTbcB+xUaZX
h1md+RT0Nv6iGOS6ZWife0h/nGUeBDqW/VQ8qGGx8qfWxHh0JJ7ZVeq5ujTNTXKB44sTAg2DiM1e
mnX/dhf+iZEBinJSFJ6JFkkItQtnd7C+iI6Y6E8oBnuoB+rqKPGDLHzC/DQlfpgwPEb6tow7NPE6
7LK6D2WjHZsNKNtO57APB7we/0ew1ykn7na9A/0VfjeNYQgxPT+/sFvHezm8fEiqcRVWgXMquLID
BDHS7cPyzm9scLQIcDdHtap3aQGxEHUW6iyFM8v2oVt2t5lCowA3qUjAL0wx/UhfofiSj1nYwDoy
2XB4sIEZnn7zJaGjbSjqwjm06St7Q/FF9mPXG4f9hekrfWJYjqbqBr+9uuY6+NdPNaN/QxFrCdVc
S4fZJhmMZc4LucqJhARx8NqKLaOXDiY6aATBg1H/3CKqIlWAx9urM9DgS+n0W8zUaRVVbte8YxnH
sT2ueUIQKFXoPYH5M6mT/FEznFPgJFsMw43ukxeiutHQ4RdjeiA0Cp75KZlTP9bwlxxq/+7lD8V8
IZYl9exh+nyF5/MVvrYWLRNBPJFmElvZr/HAklzShwPibXpaSknOiItmJ+E6nlo+r+/GYUCAaUcK
PoewH76BYr4cDGZScaMcd5Tv1+mbgXSwnH9cqr+iwwMvcp9DZQOOy+kJYbhBG98KEiJ2M6JgBdOh
W1akjRCNmBtQgR/t/KMbd3G2udpbsED/czZmnnUnKLLEeA24as6myk7jTSGQ+eYIlheUe+pxiI+6
S5tbZmuQGeje5HSGBe7UKWbGfYX4ivGswzBpxeH5L3g30Xej05j7BU31Jb9lMBgeYcIz7uNWxUum
8XeyYUzNHTJDbNld1yaScqclvL40ULCb5Z0gDbLGc7h943zAxO7+x1TllYbSvH0bWjsXB5k3Sd6M
Z30yBszma0o21NmsG7KYwzre6mss3iBUNc3hH41GBzWiQ6EPytGhozdGE3O6wh03AiGZwxfJ9iZb
0NCPd8pjW1FMZeZHcFU5jthbIIeHc7ACxCsXY8qsesxEte+pcDR8GeamoAeA4uQTRqbgiSGWEi68
dtKRl67JHMCuXc0SMnd1WKH8CFMfwn22dQ6OPu35Rhlya1HejSoKlXEQ7U3yTaLSsmPDownvv+EL
4ACEnkQeolJtWJOqIwWjneq3nwcNUl+BcKnSwtkXlnJlQZzTOMCpe2DNGYdeH1q80FJ44kc4DUvj
SFOgmrV5mXN/B8Tk1LTak6pFdp+QxNFZKQh+5TVoTrDZ7zPf7qAc0mKwNr424k3Tr0EAtpqdCggd
8eciU/5VcJjLRCv/yOq+S7sLQetvWJS3S52ylb+5F0NAG1Tq9EHCnls5NcGUelkHQAdlzHyrN27f
3s7VDiLYkMDTusfogzB+xSlAmmZfoPXkIfX1Z8hj45kjswlmB1ON2UUqZmJORbHKATeUIupGOZrN
f2I9UCv8g4ZyvGTKzw0TIH8NfkjqExJYqooRztfHTs8B93h6yLDjP173jet2R/i3Ost13ynLKD3J
0dksag/AHbV6ehg/2+kuH8tltWJRi79zHI3undRmc1lhHMEt9VVDk3rDUVGHBhKgVPaU8jcgxLWS
JgCywd7On2d+Ciav4p7zl+EX4rtYdMOeIkmUTssfa+QKuUYEvYBP5pSeherzJuejM9uNiFE0jfxg
Eznm7EmyMq0RQznRRebmxRO/u4lFOO61SKanCbMqxp3NBdfqDwLF3L6CDZYZ5SjxyvJEDozhPXpk
W86Ih0rBBHRUruvSJ8yeVQyv0Kms1O+tSc5+yGXAeYs2xga+kUAhdgDYW/DokrOvTAqJy6lB52US
6k4tZC5PtzXm+cxz2zjfUlFGg/Ds6zEjAlKNyvBmjXYEZo+anTl9SJj725UQgCGEnv9XicpRh6RW
Lut/FsJd++z49Sua+6iEKFvnrYyorJKPGXAIg/RYR7pLf0Yq6t5VkA92SrVUAe8ZNaGdSOshR4wF
iD76NtCN99Wpe6f0xBMvspcjZ9RLVeqeU3sWMNMk7omvKkp4dMRfUH3tHFEMlMa4iK+nqTV8z6ez
DnMVJW1CSdcF+1/VA62BhCT096J9NMamnyAO4WggWjTgnY2+W4CDk4Q9l5rXljEjLJ19EVbA9kX8
jkF3S8wtJ6mZfx5LTNyc6T15PFjKVxrbhaAw1Hd6aTWtJPAImkG86laRlwrU5f98ut/WXzMekI//
YIwr/qWDGnavMQ0GkOABtmfwcTgM9KZYR+lBkgmMrkuTm1go9Bp2c+dLcNvQ1QOC1qpaUlbWKFn7
rWGpCjt3FWhloMmyyBzH326wLJWUeXHowoyB/76szIZUHS3fLt53WVmdK0SZ/P0PUvUF9muZO2hz
FMLmVd4uwH6TwyhSe2A1cuui1VdomMrdvlehPnZgnx7TtUFrMiJi7/P+/0VCOvOzdvrqzVwGcrVA
cRDtdhEHarONruEuIQ5FrlJC7gAR/KFn9CafZ0uVdOoH21xX7/UND2QxYK7xxc8Y9ZksD37sL3Pq
9YJCc2yYivOO7fX80Pxug1Dc+ics2e+pU97ewcAamgxl7VG2sfg4viuLGalOhmPsICkHvGqZ6kA6
+o+dgl9MvAvcCsDu6cIpkhM8jap2b5lxtofvWD28CvacI1rG1eiNNoImz/vp/5d9/YseBJdabRpH
TaxQQUZCfjs1B5U2gVFSJKjXVVzT93S9p67b11UzQQYIAPe7HJ1rLM9yo32kxNE1o/b9TvvRnlRR
vfous9EZWTh+ucZtjbPp+CgKcPwavZ8cYsXfuMRgA/nsKIzcQpIykczJLZG5bZCYl6axuYI3ZZ/E
xRZq2ek/DhRY6QjgNcDvkV+SyfDdyzaRnAZfl2koHobCBxgV51i6YQk4V/SskE+ucBCTha8L01q8
FMg/gUmbRJEOSqWBJ0fCkrvKR1+EQ+A+GVPOgV2PhqfeCVawIE8rbTTY9geD3xYz7U+NQE6RoOJH
4PyNaw6ybTBmv8YV1Fz4zEyZ2u1SmnGAEv6+jYRKZtW0UxXXH0XJzHN6R4ZH+FDvhYHShjr3NsaO
h4/Rm2yLLMJPVVvBwWWDBeAQtz3QPadt2Q1rZd3q5bed9zfZbg3kvkXNzcCNqImJNdEgciJWAXTI
UniZQfCE/t5cDdI6TBnwTcPnjgfgjOgefRgmvjA18C6MNKu/ZS5TaJE904oLHKkMkwMypBq29JiP
JW8gjg8fqnsA4G//N8xugGJxfDEig7uNfm1onjTL6wfUflFvPoPXPivWCOeDkE5TY/zrg6hj7Gph
AN3PsQZfrVePpjzRBpG2ZLlI1RtAcALce41URWN7hnLpP1P91KLkjaLdzOt24Fxx+GLd7684WReo
OmuSuGQhpIOxCTh/acP6ah2WNH01kL9kYKAYdyeJ7mrEec+Bor7p85ealf5Vjdr/5aykGNwrFvHu
UTVimHSyggq8rLnrMdgNeeWi+zHAcXaZ4D/BDsXDTBdk1w2m2eUEvNG0zjtk/fsuMc6Lx6qVZQX+
Ksg5ZywOFts1xXAps9GwbS3Y0ggali7TJ2BUrbk4LUD6shWa97kdACkLKEFJ0yckSLuqCaAmnydc
cXt//i4twWAbDc4BJJThYdZaPBYrty0zroVZJXZQ22pnoaeOOuajjln2utZqBFXHKe/RNE8xBD/8
yAE4sB8BnQ1LTIZ0yNgz5eCqu+z+tOoE1ImFgOuoYEvkjFbFqtKockg+YP8jTMcYVko4bx0inVLJ
AAIYCFyDZsJZhm3acoZsb58p2c/nboe3/g+BAhXHwpHjqbeVrl+DRGkr2y4pfC4g2V/OuNTmBjP7
vJ0oTUpPMlghPtLUSRZD6IBDHIAWSWIaQrdZd5Y1XArraWA04Zcf5YZiEoY7TOQE5A0Z+npy1MHi
bEuuH8wnDSSKElERSXhCd20nFfXylRJAbSUrflwXMK6de0Pb+/iBLeXNLyA29AHTl0QvpLgFrZjx
+yopwVOnrE2qYnSQAA8muz5zONiPoisbJDPOypdbB3unskYb3TxfViOR+wlomr5zqPFoN16czMrw
RuO1KwLFzRoQL1/Zg+f9wYC2sti0b2eHpcvWvy7o0/0WkNU3UxJYrXfuPedz9xZavNpQs5prz+La
8GMZQMiJ0S+szKSzbvCPvlncfZcqPAExVgDQeD2ZApC8Hs1n6vBYjlPIT/0JkBjUkvVlrRDt6dVU
WnDu4MnNewvQQzapVHd7v+L7+fzhl0CjsY58COiYwZLI6eyQlj+I53miw6zRhyzwzJEacT6DSVTB
+2LlfUWbjDhvLhEQXR2BMZ5FXcZGqw0msVP/TGaxRm/fsxQ6FDs8mFlxNmrYod2Si7xOTbv9LMwv
9kTJ+DFHy+c4jCXN+Y2Ti5NoSTP/1+q5aLBtuW6p0t5e3JccWST4lnd8SJOYsRQf+Z1hE2R4Hrll
y5YxbGqPuID8S8P6cXoyij5CKAsfwjTT3ZHa6LzeWt3bsgPSuPGVcgjTW7Y3P0Fnzbv5H+OOmCXR
suQ2wR7Z4CXo9s1KIVstIK5reUpBSYV7Zesrb5k5uK6XSlY494siEXadHqPHmlGAPvwpyORxbUEg
ByipJBm/+sKsbZby+5OxvEoOlmNWqGPOeU/6f/yjD5Ruh+hYI4iSLg0K+SelJE2QqcevYAuImZ5O
xB3g59d5tVty8pmvy95Jo2glb1HINd0HROXt6923DRoO5mUL/l7Z0GQ7iOdyzNyOJucA7ZdHPD7G
nzAcbXrahXZ3y+sfgqCZHpSXDcuf8hAq6iDVN0+QD0uhwrg0FxXRUunASSST0Y1jGhsMlegLxfd9
RQtDoHeDNfGWzkNZkB5iLjJ+RwNE6EZNrE8SAG0VLqi5zka5jcUsuCwDk0ldjg3HjHOpma2mqopT
OOdTjWr3Mlb1yY4ZgojQsu4ZebpOl3v233vdfSMXWj1G9Y6gJgxOjUtLgi0buMtrk8agh2ahiIGx
CVxj1tMbnYBKx+Q21W3eCy88cwXs+oGI+72L10u4F2yVrunhUlYWFzhNvNeqaE6hxXMmF4F29uFK
7gZBGErEt4E/JKKzfkBkOVmfRJ25n1usqYdjrQsV+k71aLemoIjm4/GJAt021vw8Hd6hp73wEF4+
zNmJbIXeyyoYsRjycyw49McZXhWbHgqlWVG42uioeYYjqRJLSGUEY4nIUyEusCHV+z5nxgvueQjO
ci1tlPRpnq/7gzTiRjDld2z4KDUeJgfFZm3LMxHnqEa+HmwlJhqGhSu9Q27RJCcxBbLwKP6K8r5e
NjXUMZyZTgOt0PIXKOVH6IgvqUdL9T2rkAcOhvGyIWTVK47rDw5tLDTX6KcqAgRa6dQqmu0LhnWr
u1HQrQMRFokaq9A8JyEjGLIv5XH9N4TTe8LMdj3Ye4Wk2NFtpy4AsGwc9B3fkkNBfqnxXlvlnsGZ
ZkoejjIaYNamnVM6Q582JdDaJbyLExBN8ZOTtjFXNIAWbSQ+/1HqNrGTLJi6kDyAV6BXI4yANKeT
MXPwi3AlvgcVKEKEjiDjfX0fp2ox7jfXjRgVbiVk89LCw9uQU6p3ZMh9cKGbCcVqJ+v3ifVkaXjF
gvEIEsyTo3hmcbkAE/RXe+DccygdFNzjFn4sF7vr8OSwB/bqiIrMJp2uqnbFTyGzdgsloNPj85IY
AS1uDuCbzLJu0T4xNfaXFDsJDpYKa8fRgyFEIwNhjqDFVIN503eBI3MeO7jzilk23kT5R6ghIiDL
I3bLSHdReaW3NQf5WgoCXoCQbCWS/BK68iyibfxGfiw+8SO3bWpqVV9tQ/8cYm1T+lfCo6B45T1D
KGSql0DeHWVSE9IixOdTG/jm6neP4mML/aJj/MoiHk4qQp/ByFeVg0oG2IkMbwvxUj9bEApsYFzM
fSEP4o9Abu2fgeZtTc3Tb61Iflp9ka02WaTyNYzUbuLQAnELiwe+F2zhzjCjEe0LoCZRs617Huz1
KNCEkPzD8941bJ/KL6UE37/MYrsv9bcmRbHSJHwKkojAGf5yGgKHZGAP6hoa+fh1IB0/ZxUZVVCU
zYpxLJa8TfNiSU/AgQIeGQs7z4hXDvLG8EH6LjdBtK/H2A19WRwee9RdQIKm5yZkG8OktkB4M6fW
0AnVXoJ5TbCQIjpDUyfZy8FQwTkkClO6oL1wAytr+u3G1JKsfXcsP4e+MwFveGNLqqEJuG9I7Ofu
qvXevVS+tOl4R4QIZlMY/HvXGl6feWXOzk8083FxKoQifeThVXCYsOMXDgA9/4/3EF13IdsRSGD4
6QWd4Gb1OEch5O1XkO8coRMct0+tZZ1Kw7zXwkpzgmDgHQdEnmR7OgvRZ18R1hLfICldaU06ytYl
JMllaDgwhPBfoX2AenP4xsIx6MoV9WroeJ+oI2O31buqpMSsnNAypI4EgdLxX5NHp0kEHv3oe3bV
/8CZkcb5dhWcSawK2ii/5fuNrdZlfcMHub3LJXknSdb2Ww2Na+0ayPTE3eW3r11hIbw723GsH43r
e2dBI5d0EaWvmuFB9Ee31CxMjbYVDL1cfwF1m04HpgVxQYcEgmuiZd9X0H5N0sGQANDfvFC98F+3
HJc1ebBlpnnlWtA4eScq2y8z/Io1Zrlg68oxtQuCklKukSnwvhL3c3+/08skJbvy7ywvha6gCDz4
mEt7h0yBzsVLTystqml5DrRJZ3qCiJf34m8mwEQiHTPTyzB+Mm+rCZMEgh9kChrFVQWnqj5gU9y0
V72nCBdNwQe1KSMQKobLORPUEXsrveELXPFbwsUOUiD7P57C+9A7ZmectDJ4IHOaY1Ls74haFw5g
tlzlQyZfED5V/VeiS92zVAIssbW6aTUyZnu5j2jxwgP5bX5zgvBnSgv8+O8w/AabgJpHwdxnUpNw
ng3ghWLcdNSptpD9CoBre/O5kjF5L+QZpX41UpG3Y73AvhCA9Dw4BK+xjqs91Cn5CaDdNeNSrfe5
LGXoaffDlh6CT9iznOF2MShkWvty419v8WP/sz/0LMoygsUeW4fMvOm1fIz5Yp/igEsoAg0IoJ7+
JE/k3lR/pjyAn93JYj13cLK/+Q6VC9kVap9IT8z0VF6HSm1zRPRkiZP5yQJt9gnsoBpKwzXhztWV
bn1GWIZS8OaVNbkSKASw2V5lKoQE6IQU9kyFoaGQ15ZawuUjKPAqNA+fTaysZeGJKZ3N9mujt8lw
21gd7aFqKdDX0itJJfplySzgav/o7+k2iMrXKfJOpJu57WrV0p009lHbpCIKM/CQaBypK4BHNb0t
Q3jkvoW4egZnbui6DrQ1lPSnL78uo2BwdKyvivMq14ZogNgMoRO1LE1XGJo29tOo0rtU0Bhh3Q2u
pUxfGf9a/uh+Lzc4Q+raOHSLCDa7JeRpnY7fZIxQftwfAC13h0mK18e0VBoJhALWLUJWW3bd9vdk
4aNGj4itMSUy2zdS0EDlcTUzZ+kW7dSWJq5bqW+ngTZK94Y6piAgE+UM4qp3EJVDDgcNSkQrOVmN
Y4ai8rMsmu7/ZEKZFxWWl1dR2q5WDLmZIqYEpJQ/vvm2tzfv+1BtMrYg5ddK3MOA6q4kcuaJeGRN
af9WfgEO+L4bqqcFLYKrYGxjhfy3HNFK3KJ+Yru9tANv5UkioqyRSnP12ezYxmkcl+nTtxKfjvnu
0csCpohjwIenZ/3b+FbSH7iwVMqY3UlyCPlCpA6lzywW9PApWWCOkeC4xxNe56bV2hcFkXMsiqMM
JePhAWO7GImEZcUwJqpftwuFQamVjcft0/y2KbD8gaYThQPDo1c9zRguek//cG0nGOQM3QrMOpwo
w2Sjj9kvlfuKPjBLoUHfBekjnqkF7MsokGbRFjEgiBKN09xEhmJ2mSkcRXhC9tvVYjCzTP8QRuPW
8nGgNAJYtgwQ9G3tNoiLJko+Bdp7LB9PK1pR4VFz6ltlW67UoiQIkXvmjdBo/Q7wmeSMab1lSk69
EvwU7luX+PYL/2DpPC6jyIFpLk32ry9rVz3yG0vEof/n8YrmtViuox8IwtBizOCpX09NgMtDNU+e
g7F4Um9PKkOOqHvSjAXhdwXs1JK9Ry321ybTYDsp8WtkXJlnO3/HTf5bx9QPiQm5nr4nhIqM9PAZ
SOOaVBpTS201AISuQqMsL/DaJYWIEERCp7uK+mpKpAvjQoYVnVkuOzmUtC80ztOH1GSsbdmRVh85
tODhd35zf4ytB2mIfZNfYLSwzq9PhT3meW1Q+luxiQyPA16q0ztrqDT4vKMMnMGbAQDi/hB/T1S0
UtO69Py7OOwhUQpWJuQD16Y75VD7BtcQLGD9YknUZQj9ZeYHDIW/YiWA/uM2GY8pxYXM3v8pDsRW
LzW4I6RrI72LxU2jwuB5fjwHb1HbSeP4CBmUqMpxesxHFlvx/WSzoJy8pcPob9Zbd15rduZSkRFq
YE/jLDcyfiycifbXsMr7KZjz1XOYTZaQ7+FjE3lojP5LZJT91aAMLI3gnfYF/U2++Koy5w/y5wcQ
9mWRxqowY566Lbhhdte/mnr5y4+cfH8+WRe/HpKNgmhDOvr7/tsHXThdKDatt+tEZy5e6DFiv4oX
IGlevPeM54sAmdbuYgk+DKAuxnudkCHYuLH4FoObWZAh53DAf6BGep0glPKom1YF7X8kgZVISxK6
peHXKMI3ygNIEyCwN7fZ47+9ZB4A2zsuIkP8X+pJklCToI4YagJIYF/6Sr8ggiiaAeWdys8JUAcO
iY6rLAdgBGm4A0BGtKeX6Bxvfa4AJTPZDgk2rG8w+96JFOb6NqqAWCNkqShLNFR6oi71sxLkVsm/
TkFthxtO7WajR3owjcXddGUdF3ewC3z96gu0uxDl4scIIV8iuqDVaCCyUwsVGxVCjDWGpbcU0PQj
G+0/Ic5JoH/i6s6sUPZCrWGz9pWui7OlGmBjWoPSOQHt0nyUQJEYqKU/m1Q2gePIimdkmWzKXky8
opnufQnC9qW2UD2tgT4+bcpQn54Ok6R/FIK4PXv6xFSFgmOKSZyZJF7723NoXJw0M8fIl/VpHpTV
OaVQhS0gnRuk5tTp7kzpP0VWykDNvIlzPiEtyNSjSX98d+3jSd2eKarCZ6ExAjtZScr9YU51YVoo
iAp3BffetfNlI0ZbeKVjnMjF5IphVTxPH3kr32iWtNICrqYpnsh+bhQVZcwt9jhv5iztvdp9wv4e
ZcKjgbhBrLI6tXqSaC9XOIcAGDg0Md4oajj2ss2KFGtBXFqOxLENy6EFhvU+TbUB+7oU+zh5nAc0
1GuFgPo8JRCGMz2k0dRB/sZhA6MJmBUkBgxDMB3YT94T1T/dd+RmNZ1Skz/vnhayHM87WCv0KxCC
aHnKz/WFYXy0VHDNwGPk3j7cIb4T7wr9WbCiYTM+33kjSvW3aDlwfspMb7n3vkqAfTjfyFE85gHy
d4hyUgkD46eASiL3uEQgcBgxDJR4BtZNAemy4EeSHP1FEWRf8q1IZC76/xbuA0M6dX6eMa+lDN7K
2H+SAz9psD7JQd2cKpT5cd0UV17CfdahHk1nBwA85K+FvOLEpnxd9ULSu2SiQaOySbWqFu3Wj+9P
yGv1HaXPjGrMGFn0bDbuZHe6hE0cJm6706XLNn9620jFclXKgHbj8154EfTLdzIBKhHd6jVYkyWk
rtuK/yI88UOAWuH02p+LXDzin4bBvY25ubxU4U/XChQh8KovEjg5DhTu7Q/fMW2WdflibHkQMgzf
CMCEYTBJUYozPTKYRFLNtCnSTr767IcYRBHyCkQbLO8Ax80KCFcozAfPQYBZBxC2VvzSqP4+08zX
+2O5dmGypZML6N9wzUJ5oy/SQyEZrJuURxg2b0bDb7b+H1+sVstKBpvVn24Lls/rO1PyyG19NQTF
aPMgTQQesIFd8FMWe3gEJuvTGS+9u9GQfF1gi8EXSkxDKRF28A2GsqKsBi4zd2HOWgw0ZsOWpGpB
BVHD0WlCcMfv8jdrF7OMShcEcI+MgyjPC22ULQus/bMkFkuDetHe+PU/ZBlsx+/z30wPTLyxSNvd
6nmmJjrWgc9TZeUAlJ2WNpKCq/6HNCS343t/IIOZ0G8MrQEs9P0mYCVXymad9bj/H73M416LirkW
wIAmSiWZ39tNfJknXSLucLe96JrML/hsagE46nmK3sOMo9itUWdjXj4MVpYUbkXh2N6NwBSvoVaV
+RRDuJUadoa6EsrRXGEv0JAVZ9r9U33NzWlEH5hClWPLVsal9krPLZaraIhDvbakfs50Ivt33WJ4
bvBNRMjhKQuMTNtvRgQwSd8dOW4sNFjXKaLYzjyxJX5sRdt4W2AOgiryFp74mQEnZnp9uqTiDwg9
MpFs+y4mRCJPjERKZQ9COOi9KMiQWdTdEwZEsytqnWsfv0F3e5vsbxkDUz4op5VS7R37TpGNmaSk
oz9IY3SY/7ot6YxJa0ni4ZF0GGQszPQ+vZGZ6+mMShpURA1muSVRD2mSxdizHjlA/Yw4DysZ37y2
4GcILMwR07YQXj21idmgsTmkF1bV9EDCQNhIUdmDDyvgNoXyhCc+cbJBqPGbqI8IFLzy/nq53zhP
bl8zxp1yoigpSPSMBFAFKnYMHM63lTygu8Vs+uHctOVr9KRMN2ZMxxSuXqgoZOqCUBpUct5AM+zt
k6d/qMhNkv46kQCpGoakFVP2s+9kYjrZ7LqwffJoFdeyRVV7jLNuFOdY59T8mwN9yy5ZUY4t4YVq
bo6ZLXFjjvge4TMe3Pu1wUxtNFGb24wbSvGz7adkM4KVLfyfyAnE4dpeo92SELNdmxBtf6KWZOng
zQ9dAYTpFTUlYIzIqFHHL0W12tNTffrMG9bAwYsbIelMzKTqwHZob6Qenq7SPQ16MEOpcBvZ5eu9
s0BUWR9iDSgC0hlFNzXfptPT+O8LvSxvWAjrac1mnm0ngsD1i3ZyFsssUnqE9GxIKdEbOau3uKQX
BRziBKsOEAuMLRGFKOUugJniaT0jz3YVvraQZcxdzVe8dzIWGUbxQ/7mtuRDCxhOlaRaLS6qL9J2
DsD1Bl6F5yRwyH4OldQ2kbIugX7qTrfcTLlUsb14PhHEv16SzxWjjByJ+b5ouQ2p5cYXvyrCz7Q0
M73sASYPfAwhDndOBZKCU1ds7zj9RhNUMK5fvlWYY+i76O8LqwC21fmHqg3YTTY0hQ2oGt5BVlcd
Dv+awmukZDvzom9jxYwHAnkSlBVkpWln8oL5zVg6DPu2+3iMg5dMctmu4ERC99a2guc7ksobbtN2
wzTtL+IyevzZ6BxnX6ueICxNxmr3zdsLNcIIRmj0QstcMSSqPhSls7f/abB2Lb8wHbzEOtee/mV5
Km2SoNYtc+mxnSVG67xu2ChPw9DnohWzZIvrcHPd9manXxmBFInkxF9H9OTOzd9WGWGWUQosrdcK
1fZkt13mGCwwlFzfBk27lvne9yhAi/Pud2GtS0tGcQBDTJkB4wk5+5knAjrsNpszNE8ieOWuJ1Ym
LKlLLcKGWvTvcvoqr4qOpVHe4FgkqqyT2OEC39jRSIv8RqQ5Izpm6kYyDUWn/8OHC8xhbpT256yl
9vaV1aazVOliFdm5rCIp0NtFFFR9Gv3w3tAGtB6WplZp9SGduhF3fG81vyGsM/zuXYMGQNl48nVa
QUNIeik+qLr8Qt1RXgLnJGCYQtRd5bb/fCSQ54o7eSIeRHaWAZzFSA9SlmOaWk+48xpeAYX+B+QP
qANpl5ebeM+ZG3R0Vr064WNRdfNeIB0ODe6Q6ter9VOekbpbABXoKUfDlmE+xgIOAN2DC8KqetkZ
q6KH0r5nS0SPcNePSh60KBGQq57RTxuGk24MWMV7mtNkXGkD8+gQZt0k2a70EAc7zkif5nWiZNfw
SFT0kwlHpbIOaRYbf5hKsGo/06Tr7ihnHN1UNwaaNwPKnGtAZDyuSj+E4yIdALuD52x+qCdQzq1f
WMnyRTIjFUBjNpvrdrX9WzWT+2NkeTMyNn5F6jPmP0t8uqJVNl1HWBXpx8FhonEjQyg6DUxGrp9o
aZq1D2zGf/L3H1D8hg3lt0LnWd9vBMnEwy7OskyMqZao3ZiDrMZBWeAzXhuKF+B7E5uUjCws+yFW
uMGTXJWoXWL/tKTAtBwnmLx3ThV/ZZOVPFA5SHVYPkiJJKFqehV+OX8SWuXDv3kbdj/RkjHoRUmu
qBoCDxJUE7LQI19TmQcDOQQ4Yys/7426wMw7mkLPNOBwFdICbMzhow5J3yQJy9QDlsQLH2VhK/F+
UE9WXE1FVZnQkrHsgR3fcigXpF3wbqIcAcVOSE+OG1CgAVyw8HbuyfVwPduWMxlMQGmDEitbWRyq
RfQeIrMbLpt6uyN6gEXWxPOIEUN9Il1kN+lhmOwf6auvKuNZ347TvNF7UWWYuQdPHZujh+ZERt2l
6DbdH+P4udIoebxfLc2wWgI040e19ICMyfQaoDMi9SiwRFAyYeoDTo8wetMze1kelay/1Wvvsj+F
hj/xR7FnMSDDj0/N1rUsCFha2dj3FiO9zgdIcPZixKrVAmjZMANjxTUxpcFXM6ROxvK+7ucpgiDn
X25YcIZfgqRVJbKk2WOxFI56r4b8sah84ENTUJmKBrs3XJdbVzfwhLetd2PtN9hm+qOJ7LUauZIK
/OjSa0KwW4s2VFQUCEmMSEpRi2a8YFYziB4OJ26HGhnq5esFjoNebLkSbHBfXXh4LAqvUQZAecsj
N4IscZcO+miFPGzc4+W2JxJ4jXqMZcaJ/gYMSCfLNSYQRYEsBBh2Lhnlkvln2iNsnaasBMor7yTe
wORPCdKVgrOIb+2NMTr8S+cNd/0gnQPmfmHshBQi3bM3D1ggpnU8ZXCoPm1Qs8j1ghCFmoRnVCBV
ggCPbFa1rylOn42KZPDjdxbOoXKDqxTpmUE6l6itTk3mp/zTW3EE/QVYd5q7puB2Gyi/eRLQBrzE
WOl1+EduQ+itWtWzp5W1V2powe9+2bxsmbpLacDD2/oEpd8HG3GMc2qa2GIZkVtKXOBnWjZ2Qp83
DN9J6cGV2Cw0zc7kYRPkbwtcrNSQpXSD6RohROcqSZYY8E+leiXMtMT7nBgTA+lI6YRPFIk1hq0j
IA/CFf/NZZ/4Pr8TVaBsWcbf7pfiGccyzIsxroms/XyYUmrImCeeiryzK4S21PrvqrruSGjV7JUt
bydxxtjlxRurChy3yVzhRoR87fMqLONYWt/+aLn/j2zqKmbW6HVzYynfqf6VqfGHsXhltGGnPC0P
hE4uBZ7R1j39St+3pnpxsRp27RZ8l24agyxBi+Mdv2iQE5xlnAbNAhBTPeSB3jGDtseuiACZ5eN7
2HEid9j/XpaZ7BpS9OCKtVbwrHIIfagZhSJaDyXVk1gpuvNxreNifHYNZxj7340rdFFQpKmptKcw
2wihNBF+zvdbyl1r7D6Xq+3pulCzXkn+o5pARoby9fKvGBODtFsdhM3vbANYy0OtAzKItJVHWo87
kLo74HeCyBRvOwzCalPcLdFOo/0euLBcoarJPp6yuhV/ODGO5qnNHSNfsBCO41sqRXfHw8tkacgt
Bh2s1YeQWWs89zisWxtvvCFRMduiKv1TbGBQdIkXY8FXMSjnKfRANbRbL8xwGsA5/faTmqNCO2ur
vTgOVk+wv2FMmaOUPXThGyLLI/zXjcWigiF3UTK6VW+Z2IAblSqLzsmuklatjKelZ/1031DVqclU
clQcph6UUqtMnOsBukcOYpbN451DovLle9NgUlSkHCOkd8OpZIWmiN/vfNpC5nnpK0X0BIta/TWK
bnQ+5N5LIH1TRuSxgcu57VOlXqpnlho6n8kaq/hEVGUOCPE6hV43lr/nUzP1ZXTybmTvS/9qXUx8
SGR4aez3sXZupqy/Rm6BEhE9iZ+mRXzS9uqaMA1RY5NAKmefP0LF3CCGJHh3Pn+/CRMke+GqzB1w
VIiRvZyiQi+IqR/cPrj9zhv+Ukq8tAjsj7huGmjRLF6PgqaoZEwYMvpTm9GX5iC7KW7SG86g6osA
Do/AHQE31wWzwD3aenIKNuUMkh8jdbTtyG/gzKd9vKO21s6/dxr/qOxDFRv7yPUEbH/yorYu78Hj
uj3MKxoAtEO6aGkLia0YqltTh9Sw/M60RXxcMGo6QP4ouMRxRdZoJqBArk8gQGXT+ZA/ygC17rKc
xaLtF9PrFzy9qm6gG9nmbOdL4NgSuXO+0SUkU0FPDi8+OvmCOdxykOK5clPQ5cRIHMCeFa9+0uft
b0+O2yVHbhVBa1X0QgXO2hd2vLkEsmHUpf6jfGq29GpFDPuDSv4v8Z2vwG6FI89JrrNG4NmWXJr0
HtNPGpjVfM5u8/9ahlHtugxro87m8fjBvItpUgVXsQ4FqLXLSBCYtEypkBdKEwkM2GuWJPTVf8Ld
C2TlMAE7DD0rjXemdT83FRiJhdQXfYIIhTljYOJMomscDlqVe33l3KJfP4jwGGlPVPLTuGy37llQ
Z19T5kCeSUD03ch3YOEljijtZhtcGrni24RuNPh4LPv0F2LYFbk+iyW7J+Hv0Dl0lcQdgVJ2/l60
UpxSg/0YfMB+aE2TVJdZFXeMr39swxC2PYwKUbljzU2ynka+SqFjMjT8jbbg7Eel66VEviGMmPpn
v9i2OdlY4JB6SJ8mxEqJ0Y3hQyf7QGzBEvFhubocgV7u3JZ7zrDBmW9TpTc14mwD0tC/0M3i2wad
LO8f+YnYzdYQGrAt/6itKR8wvn/prqE9h1s1uXd9yPmRJxN+t97MSj4H88a3gGnJ93xmpmEJKTdF
JZVf3s7KS62CFJ1dcLEh7s8wcmBzruB4YStIz3mxKDl4+vdZO28jJTSjNmtU3XpyC6v6jQpY6k7h
YxzWb1O5WbvI+R0H/UNSPW7uqRo91IK7VzqXR3uC7hE7zwUkaWWeYDq53xxg/1z332LbnM4MUJDe
a0gG/wjP+F98BnxzMnIdi00M4d4HqF0bSWaKHMN3KYEBBPzkT3ZaZcRxfeR8Xelo9CPVPfUEv+h5
HmOoka2jjeMzupjHamxHGZunFq3By/yxyc3wqMK/n36k+h4XaCk4LoPXVq8hpTUXfCVpDQck2afg
lZbRtV8nZhsmxhWmWx/nmdDDvphPRDbeLJO51Jdms6VsUmfWoEPk293CbageVA7vEW2m0c6dYUNZ
6y0muy0Yl4Yt/dIxIBT18c2XTU5HlHU7VHZQJGjg+MB+CrN82iEB47Hp5/oRZmfDs8zGmCT9oHlm
8zI8eFp4IodNfvLMpCzGn6S8YEFYTww7JPJ6CKOHn4nSZAr17WEAz/XsA2aqGU4Obu0bSeHNC4wc
xpCjQm5Lgd5m+lNaXUfmFuLnbGSQtx1yHX5OHaVBIWHzZEV8f2qgr//EMGEBcHuhRmu4K0Ddo5ej
MZ5n6AMaNDvzN40IIVpF+G1JzjPQal13nrIurwYrwZSSOFSeGsI9Bxpt8nRGTGaG1U3T/unOqmr3
GZyRLdvBBZagDCxL4nVT2DtO02tnDVUrvyEmD2TOk4aGp9WyHwE7nSyEHVW6J0A8mdanYbax7lKX
Z3mVGQzQPQOya5Z4y74pWWX+VjrieUIFLfM8R/IQFa0BGEMx9+dBbWH3GcJpq5rQHWdPswtVp34E
X+M+wgWOcOkJxSXIzdkonVbjkunhab/SsQm5OAzLdb55bRVWmNXCyReqqVgqCRKXEquRlXMBGJqm
NnJIv3U9vZ6iLXwfv7y5Czxn81SVp8/WN7o4ETRT7EVyPbn1saer74gKX/lVXfQSxbkKdnqCt/qg
Zi3ehSiQ16m6u74cbixY1jD/vl0pqZOG1qkL1147bhPZPGM4tO1EmXxCoIibnRF5WYbNZbcronF7
OAdXCSqovV13+bqfvwqk1JQRFqd/EuiC0YeMDkuvnIaXiPog9pINMUPutcBjnXwSPx9jcjjkD7T0
/cjtgLa5n6ys/q5beXst4PjtVTwBfgYHPGi1vHmPBoWC+Wc4CskWE/QYq+HFjRcGb4F7F/dz/rOg
dKRiELFfWwLwExxxN05XMzaaiKevRGfM19ctFu2bNlW2TIoqbN0/NINAwBmI9B9L5zb0U62G8c2k
i3S21kwNv4ox9nxa90DAeUpfVM3oHzznxD2b5ln9M+E5qUZ3bLmqoFM5LzJ6KYYl73UDm6pNJR/h
f4kNDV1jEFiav1Nn19YIHwaEh1v5aCsH299EMN/lXB7uCENL6sJzSrx78UmEJgKgYQZ2MPQBgSLK
gItsyq/aW2eHWu+BPyFxpG5KXnCxzv9ac1kg/ws0s5ediq4FIQqhlq1/6OMYH8bMX9VQ39rq1yuv
R+QNKk7WXtYUtRWn+hubnjGSzw0kbbCp1eoEG4BjvL2aecKj9CDU+lVgZhBstPBOQiN5Cqzm+gTM
wl7KXIpCUB0hiUd1I37e7G4VwA/DBfXGJVc4rAibOHaqiR7lVXxVubmCQgZYalztUexZ5EVzIkGG
Mer956L1N2V/4w2YosPLYvdwGYMxtIthBBfgzA4oOaMBEGtHT8mgM6TwxJmryqwOvwGAPJamrKAA
p949qLPWQz2fmqLFfYgFbg+BBX0QGkJaNFc44xzvlowthmIDfxueDSbFXV8kr4ZAI/U+FixZ2Bu9
EnI/Nlvjei5mrapCz7TexOayZGR3M2lqFxXUhD1Nks7QDcSfmgm+jZo0wstJLotGyY8uifaQLTI6
bqB3QnlDZpheesBugu/pnwyB/QlSkTBECuGj2UGCmEvLHvbQh7xN92ky5K20nhNAKfNb8OHH9wlh
Na3Or5KqCk5eeytU1cTJ6AkrPNMNaeXkJZIuD7wroPvw2q0fXiKliQ7bOwa+kDNwLdBQ9Y1Hpz7G
fMtRapTAWoAvuEXiVvs3fZ9zVdM5kL4oeVmigNG96csjnkzKgG+DlXMsnSvB5JmhQ1DZQD99v/84
q/RZbcb8CvFGOFS/ssr57yQHcptSbdMbHx9f82U+VTk18QVCcOQk18Vn/iRLeqX0SCP2HJTeWX6i
VhC/RtV4OOLVcWY0QqTIZujIFITGAxBJXx/HPijjrLsjLfiUTWO/s5Kru3Lw9sSJ1drVLdAJZeHN
Kqg12rilhZCc8VM518ZtHvcJun+HxtVuQnDuctN2sHdPZAfxde8M+gTxBwqmCmD45ymedqpo8b7G
3I8R3m2s3yiSDG52AN8q4ADfE5pcVIvobjW9RAhTKp/YlQW4Gb5Wiv8u2g5hIh0+bGs6YjSvJu5r
ACzJUw7D6ODr5sinsY1ezmlYg1qRF4jzzO0j8kjZh5V/Euf6OXeipwDYjRKwbkBC6gnUIhOcP/u/
n5j1PGNdk95dX0QnSov52u4714uTIr9y5m3tDq5t810sLYs+Hae+I3NhDg2c2tWpHGiAfkCqsolO
S8LYt+U8VNpuG4MDvHji0YPv5U0pHo1QgwqIukoHriSpfs4V0Q14XUMQBy5AXySkOoHnaIa17Lgd
Eb4ZlbxUEizpOwkf8rGbXeRXIZlkbIqIYsrAml597EPoO+ivOfbDH2l50hosc59wNIPyRBo1xF3g
+gA4LWO8VGMavlJ76iWCuhbaK5hIRVfId3iU6ptjIan3prGWQMjAhIYkp/uHYkkRqwIp5CDLbWIp
wS531W//hXFCbFU4YLEEuzGaZN4jj7nEm8cPmV/t7HeOzTUrxD09PZ3ckRGb8/xTtEd0YrzdVaLs
+GHIX/HIRmW1tgerkcTjAEMT8dEB0wS8flu1kFWvSQWAKcE4rBfJYfTEHSGEucqnqfJf9GIAJtg4
YIHeNGc/YIk8RjfwYtSpzKSbgyBOw3TaS52AY6cAvICmaMqAHbJOUIFgqF3btLoXlQOUEms85rCH
r7V1qcEcrh5VamZ5owLEeJ/Mw/1Pxh+k7nKnwxWJGW1hQ88yJjGJfd9PwGwBdVqzQPPMN+9i0QEU
GqsKrvVuYHcjzuATRmkm4k7Y9CBRAVaLkb20T5A0XhXyB7IGZEUiW7+guSp2ws2v+OHtkCxqmCwJ
vAx4BctRhNgKC1JleLdIbqbtMXrqcock2w9XwlGz8PKbrlMPYWyRxoMnxa1t0V64r/VGN5V1YY4p
JxsVtHwtpiPw5FGFqcPFdoABrZM2/Xch41qET66IPgzrQdgGql9mDiGoBw9fDW8ptEQlp9eKYCLC
WzXS99yF6223PqH4/ymMs9MOiYmg9U3EiU0wje+kbHxZJvG5N//hcAAO+DO+F3Gi4TTqAyjlivjj
qyPki4ooQw0UwPF1wdrWbc8fjtaqjJIGUCpxFLfRRW+7sCt1xINXFGcZ9B3XuXUV4nNIcgvRO5I8
Ne3LO8NjcpRp8AUzFReGgD45Z5cGqM8osStENSZv6c/6wAwxRfONJplqz6jm+BPCD44Ve58PyEfD
ftdc8y7weo/H8IqvKe3T5U7+SvGjtu5NGxqu8NHsfGynG+mAc8E5Er5wDu0z6zujpGDetkxBIqcP
aKvVrM2HqMKgwjda43/nhPiBqYmXImq6OlKq95nT9ri6t5ZsMgZWP+OGRxgzR94g72wj/EoKOPJb
mhSBDp6ui3B+PrqzAFQKtYGZuy8672KaoKDmXzAv5Prf8Bj95iXDltoo31VGleIG+de+GVqz6iza
y8O7vWFgO30l/fyBpM/CWdKRVMEjbHr5LHsa460Aue+8JDjhR/JdgBuzE3xSLzSQ3qa4yHLMyYyU
vPSCSflH6r3uwDBobQEJ79snM0JU3fKg6UmiKhgfjrnm+Rg6owiTt4lUYgkHRwZQlCX3jMNtnOlj
YVAWwJvhP/ufXazXF3drJb+aDxJizkmyWxbsXOi1o8HbhEhBtWsayg/WBddSo/3NAVdDLhNACXeJ
G/rNiOECUUWVJCVpnbmVYOYaNHYdUCTJ0J7GltXwH7VOGG92f96ewoK7EtRA04P7kxkQTeVYDAq/
Yj+MxTpXANFR1h3lZoAhyOhhqWtJqL8rlT1JdMLlvj5YjFy5oPlHHxH39P3Jw2Sdsrs0Isl7xmrC
iHzB6iFOdvlaymfQ/PBqVu+3LeNEM+ssqrqyis4edYS/Ij+EwZJwLY8LxwrxJrjISdt0GBmy8tGD
AFqIu4QZ4icNE8bZDIuf+6Ojl2+eWQT4HOEsHkIVj23kXajmFATQ4jyCqkslhqMjfNi5H/SnVAU7
tVEF13PqJ+x2QqOwQ62WVPchFCI3J5dhOlEcUE2QTGsky95NkBSNOtEEbwwBIi9kaPOm2HdLKjyL
2y3PAHqY/d1HRmxUCSKc261RNR1313FPkmja4V/wkyjNzO5cnu42WbqdYtwFOr7PgXLR2RYTfEGr
2pSBZjw7Kr4wLaqwkCt1diJ70hXwkrfcozZBmBfc31osrfOuqupVRLNxUeIENA27R+l61SQEwz5G
v3dFaOtp3dU0Yr2gcPxZsgRi4uY8Pai8VzfqGEHHIO7KzLOOEN7JXxl3zUBfFYJKZsoeBMRFXoun
2y8cHWPZl+bZrMu6ddvFvMNnJ3Rxc2Od14RPUF8JFiG9ArDi3NLuOnMrOBDgYzaGguTL00vESvLG
1nGBvpO3/Bn/EzbUA5hWoqGQ3A5O81FXGs1LobvgzJrvT5pDw2tGerIf3ZZYl23NmqyhlxfGGTm5
35BnWKcgwr3X074g6K1ADP0UMvScaveBNOPgfvpZx5fqQm7GB3Ohq5b3fhz6D6B1HC5qo2VFIejh
++0RIcAkOZRmMukxf25FosuqWZan+1RHdtsm19RS8BxDl/ehf4pp7aQxotZJG3fMIpdl830aaRxV
XYv3sk8FSuK6In2PlKgj4TLtrujFKdC99GLYqHHUTUBzqwKudnBDK+VGE0qDGq5taQam4oPp20Sc
NU13pccvAXCDPNc/pAKov1vzI/MDuzuGc1csciejjQFrPNLecAEsOzccO049GmrQ9519kmRCDm5q
oHQAc8OzykfmHGZ9E4vGtOiEq5fSz30t768lvnTMxSYZulibKSCoQhMX2mhMVCHD0So5RBHWTTS1
iHj7i06CvAeWmqYcrXMG1QSIh2GhjBs6cFJNVeyiqfzZO6JWFvxJWeXWNZnf27/rJhvsRp/LeZGV
p4ASYBN7Xr3jZjjdSrBQr7gmFs7p3I7LNYlKM2ZEoaOul8Bao7C6ixvolIgGLLpDBpBnKrEBaVjM
gW9O5r8/3b59mom+fs3Ik+Hb0ZsDuc0jVhP2xYvv4whhkuStI5f9hzLP75jYiMH755clH369GrU4
M2qXkDnhn3ZlZryTE+C+G32s1DfJ8v7gmZo85RbJMy0/PjVaHkcQPruFvUDP5ICeJYnXIAvz1uQU
Oe4OBi26hPEA0z+zhFZDRxNluGsPhKVhEG4SHJyHg9N7fno7iyLBOjlMP/sT9KbNZOnaq39Pgv65
hpesVw2fsKHIhp1QnNCEvnil9yoAIcLCSydOK2rKVX2kPyyKWCPlni03dz+oTIc9xuI4YtfCs8po
c2plziKkaqzc7XW6v/hbO01zhU6Ms2Ds1zQ4QJdqJuTHwAIY/10+jUM9xQSjMElWh28nIHyC5PEu
CKwhHp48ZjRs4Rm7A8zfM3nb4hMQF9WUi6fqu2c8zJmOXJgzTVWdKqUWmSWi08dNcMUf1uiM957D
3VbEbitL5g7WQZ3M/kCVjbP63y1oYcHX9n56QACTlepLpSMgdSdBizFLEXmXrcp4TaD2RO0sRvKh
toInAVDPs84VNp/43Uw1YSfF6gc3W1KSleLwwBxES3nmaLl2Pu7t6m2vANnR1XXjFk69fprNGX8C
LkgVDowzsqmYaB05/gfdqWK0xggP6Atn904XOoPoD8mWMSAEHmkROvqAsLGxYOX7V3zfFxzd+rqf
EIXeCGQUUaKXzpnN1D2kMygdAAcTdbYmJ4H5yHLjGmREYLhpc2DuEqJR/w6iTnbkPY+zfdhJb8J2
KiVfcsLf/DpXXcAovEvqfRY1ptW/OY45FWtBwc2eP2poH1l/qZ7Dt0992xxpDIxWxCzHdppfzpxc
hgL/4po2TxWQKPemL3qow9Jo0u9dmFSIpXw44HIHlvIYywDlqpgiXqHUq3QoDQPe/NwguhpiY75T
Zmyk2qyb0H0TvKN3g+KUmqU1p6Ta+0c4b20FQdGZINQJivRn6fcxkd4qqXWqQ8bLC3tZCxvfb2vc
6dq1UJXpLcF1dnw1lvK7DtsUMZUuxsTz6dXrBl3QTcKGJbuHC2BZTW6+jQKC7tGh2vif8LQjbwIt
UKOG5mE1+FCkwyb7A73d1ByvyV0kTV3579hUwF8vjmlcrw+ekqGpKeLTaIF2BUTZQUGtpEuL0reP
H47G0jw3BVlFZT2REseGcxs43HpvzKuMr74EZ5omIhTuwdiET3cAjQ8YKj7WiFvgVBmYIGKLwRO8
qMb0RKjSPzRjvHdPt4o9SoGQ996bKc4WHr6vNFG385ZTiHWoDqvVNsnT5XhpdCku0Ur3vwOaGCEf
ojDW6H+AWNUMrW7douPHcd1Y4Y5zXm9UAy02LPZTbUbhygn/NNwF9DqL98JUwsYi/1jUEvAMsNc8
JerQQgRC/wBUBW5AeQty/iJmpbitzyo40mPdaYO0pvjnrwsqBWIgGD85T72lSnrFD+49nPRCyMm0
AnhXuxtz5MpQLu/Pr4XIidDgDv44VkGbGZZHB+r3+VYz4+eEqrM2e1DooQUryWXaIZox6UxA7l4i
GZIoqFL3zP6t+XtlbUpTOpgKs7s9qhm4sC6/Is31KmlHHBjPn0UFf4NZhxM7nrCw8LH9WBAAlonE
ODBPmI4brtynEg+Xx8dMzWyvZ/4JJC2Ig00IaVC1jC5Fuesu0l9AEnSk7BUEur+xo5W5C59rrjY9
KETjzRclqSHnZK3eIOHNdc0zR9BqPAkZCQhT1MJS0TUrBExjh3y4vKyjoy/8cuTlmA0LLBJeMFO5
4IzcF31c2zENdB6p2U3n+LCn3XjMPC3i3+nF0NHD+dHg2ZMkyvM5tSpzUMsbfOoYlLpw88TLKFBd
Tq5q8P/T7fV2c5Obrd5z/IkkFC0apiQ/U1Ub+UMTLQXlB2ma9sLEy34XDsItkSDEcN9FI6+yQXm5
PoV0I0ym+CYce+Dz19LFzqYnsGXqfjJLJkhdhU1BCrKeJBJt+FFlQ2YTFIFd/yTFveZMoqNpQ2sf
EKpYVa4zHFieplaKQkErT0+vrfmP4ZIsu1byaDCX59aX1C9YMVevX59giA7AYuyjAIIelShe8S8j
I/JMD6iJm3+FIsHgc4WlbkPNAvbR3SXJgUTGtPcHKdSLp6wiSsKe14KoFszRoGgXR9dzPFo05+J/
TpOYoUaM3xznJCUi2/wIUv96A5x8aIBWXZDzj1WWf2pHCahZJZxJXf2puoXRFtWvL8hQH2tDXI/t
16bcuA7+uw4duEN7mYBsg++xTumBTxaq+bveqidwWeX/FB55xYOGE0/dBSNWHGOrrx7WrxjW6ytj
zJfJdbYrK53VlibY5pvzjU6wayZCO8x4rb47owx1R4qdR8xE8bAUy2KuRskimLmZaY9TlaLBuoVP
TeKgEPcwtZ2O+usDADtYGbkh7zZFpL4BYXCsp/C31TuovDutKTMxnsoiY8IwWK12paeY+3+ODfOQ
yXANu2z3FzrRPzYfwRO+wExqI5XVHakNdzpif+kX4CJQIhY+Y/0fx7gitR+HAVooQtBWRG6lqGBd
0JjzFGXzQnNHJGoAHBxhFXTGAvYJrSD+Y79hNO8QGbAT9ezpvOejof1tq3jPoNUdQBscGQ/0LQvM
jEoaHwVYWVqU61AisDEQYiVrIeamygHbqZSHGZTX7qcELNE7CovgAD0xx0MJUULjOnqfCX9bt9vY
9+k6F5zOoxJ1qkq5LzAq9kNpLOayR2ysDh9U8nhYVWl8AouQw1HbtLam0wcpd4bq+ruBraxne/LF
f25nt8pYLUJMb/cib2oJ3YN8/VfF49YN9YXSkELWTnG5nvs18Swufdot2IjhdUbrjX1JslrAUe4l
NHQRZqpJXrHt72AGLrMyosnuB/BvSChb/yh5HFRr4CJaU2UplALMo/nboXwOlUAEMBb9Txx2Ig1a
yTKaCT7+kbhC5oUSikYltmvTip81K6Y4/1/NWSYJTmDVPgzyKGJu6uAbed6tCYS/tSBK+7Y/ckDt
fplS+ppQuvmHQKE6vseqvXyRFxG28nsw+RnL73kCRtmbOWPSCSWm9dPtDqIZsC4447uhUD4GTzd7
z9bAnuFJ4eUZdhmw0/fhI5uJBuHeOr0k+X2t9ptVwrGlcWeF1l5EhsMpLo/RwWOmP30UhFX0dd15
m4Uk94Sb4cu0zeqqPEri8uJCe4gwcvT0EFs9pu759woozqNOg1pwZyTCLH18FItTg5C4uGERVWtK
z4jRqaC/DSF0Iv/5rT9ll7EHebETf+joih6k3jflSPBVQemivlR2rT24y1rJbWshtVcp1PGwQZJK
i6sMGYIiCYK5ravsIZJQT7BZjt9/+AntEqjj6pceZcGHMuQj/roBQ+jzY/YUmRkV8xoERFGtXlpQ
qfDR48StDJhrJJKjXnwjf2my0a2clCMsUoYOWPGAogGKcUa+7i01jLlb0+pwrN5sz/a+tZr5xfW+
ECYHLlGChSAjQeUh6qGkizNxqDGANQhod65zdLGsB9tqD4vsTdTdxP2Dh5GtGjIchzYeKuyPu1Bo
QrMYl70jUXMwI4YEQ0h2OMyX9HwjiSqSHG+qP7SDy8AO/Pguor01wMLBgHsXubA93iv/GPwgqP/Z
9pmaNE6oHTjQxaJfixJXbqslBrODTLvOh3PRFroeOzWVjHXr/NCt2AfrpamHOLbPqrHA5IIbJMT6
SZGKPFtP78OTQbtT78+IoRLGWIEFvYvB/khzHjuYkBjO+LswSaynJ9ubKphOqswR6/JXWRsmNdV5
Zk9kQWxFXXRls8cx0/KVjK3f7WPqjb36N7cpLr0dEaE6Grzj4BJpjsGRDQNW97J5rnCum6SvpXV7
zLIoLJqRpaYfrkjjccAUuDoIowdhYrfCnkNtSohuGyUUfbHn3VQzOrznaNCOAKUVGZ/7RgONiAlH
bo6koLEfZFXUfvEOEZSvlepbYhLsYdt1L9VPKcZqfRSm/dFpudpEPLg46Hr0hIrlA5DIZkUS7QQU
j5VIjszB5G5eIKA4Geol6AxfF4VYCm5vnH0OG6jT+hJQmZ3Krjclj4Q+jY435Fxa7IRGJiAUMNfK
LOgaPZVawroj2O87OIk9z+xKG/8djH86dSeqpmuLWHI6H1mlHEXKDXM3viNHrOc1/I3gx1Eg54sY
xCS2edhaoFbB4YeSpY69F704OPAh5htSofxfJP8Wmvt5Yqvv6mwCAVa5zhsqPJBKN1ojzj6iKNS1
SfWI8MZA7z1jI1owPb2nI1Bz9PQJFUV00AIu4euQxbocMGK5uWXQsf9H8oDGJard+aDqgd1XdM9r
gGrMBDa6jaD2aQUnj+PPFkozZBzl6OCQBrv26SCdnPDqxkNsV95H/fYpgjj4M2lCe8BvBSYKYxLs
yJ7il71caQG1Blc1zpDy/Yax4JQq8WC/Zd+HbtMyPtjm4Nw0QnhS5jqytQzKuXrDAEWFWBjzwu0a
BkFV/CjshfzdfEIRcs8dXH6PTJbVGKyn9F5SG94sakzeG1Yv7YNTYYwDmk23Gx58kZT3w8j2D9qW
BAe/hXn4UKbKccgg6C+IjVYgldkbOR71Td1HYbQqB1JsQvv4stJf5SeG+83EEuYxmVFwgAbpIMA6
fIjxTiyaIezacAFMwLVJN1Dne32WIVRUuHWSV+VokBNtU3tsIn0KLCjRS0QjSWrMppdhFS1auDMo
aqKuxn3t+sdmPLP2m00MDwN2ooJ6wp+qr3RNi77HJaWqYWNHuPLuCZ88hMLQAbq7AZlwxCJVLiMv
jfVMqprcDJp9v5hsjbzXFPufruilnIX5QEW+emzFOJKC0wYDHmwIlJ3X+EMAsa3yHeWbo0borKD1
mSwiX7yEqWkOAKFHtka3wDXz5oRpLogb0Sk/aUTeCDnIIzNBhfzs3OMq8CNt6eKdRHgjFaSmqUCJ
lObKYmrksBlo87DYVitPNPpMl9XJQKn1pj6QTNQf7NEgQOfnBS9Wp9evY8Mu+Gzu1UWhfTqNO5HJ
LGPfJxnVr3fE0TPeEU7z9Rkp1bQ3BQH70C76QlkYCly+YC5NK1VBbLuHnL1oieqVoI69whRb6URz
I2KMwzlLOK1iqxadiqD7KfpN6TkzkyjOn75+tkpyTFDFqL2FcNBPUIQTg34xNdvAPNN5mYi0VmC1
BVXS0AnuYMVSRFGAf0Hvp9fSN/Xjxc17X9DO8sqKpJsEIf4F0Pcm02yOoJgkfcuoXc7R7dfq9m4+
pHC+6imHbaGlcILeh/z5PEfdDa15Eg==
`protect end_protected
