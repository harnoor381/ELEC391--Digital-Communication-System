��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����,�1	�)��&��(��H����dP7ɨ���:��0����,�6m���Ib� ��JK�yUh^��9���E`���K�
��Q/��V��T�"���-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_d
�t!���N�S��گ/�TNM{�C�5���M��;����L�S�:�{���\p<��)�0W��B�R<Qt��Ԁj,3Ӂ�v��`s�HW��眣�U�Z.͓k���ŏ�^�sGt��P3U����ŷ��T'�;�5X�ոp�XH�>/_t��j��9,����T�	�u�M.TE�hV*���D8��My�U�z�$kZRn��U�2��WlcgF�Kd��8iF���`��7i�{��3ڽD�:K���U�����tpyY]V�*'� (�u:���������!�Z]�<��W��0TW�2cŹp�l}XSH�|Kl���ԟe����#Z=	������ŏoԻ�ߢ[������!�U%��s�dO�����_H�4Q�3ũ1���q:�oͲ�az!�n��i�l{�	h!�r�g�(���;�[�YkoP:���4�_�mY�5���u�cdԅbPW���,��
N�����#9�w�6�cO6\{�ݎ�M��7FB�gt:�	�R��j�i����nn�<y`�N�&��_��a��w
�1,r�N/�LOI�k��x��Г�����4�K�M��2 ��rt�`�IL����qza`�4�n����g&���	��u޺�Z������k���+Zs�BXP�]=1a����y(��5�`]L��=L�� hL�p�{n�C
�+^K��C|���ʻ˿IG�eci���,0K���AaM����t����;e�v�4�j��si�E�gh�l6��xI��)�ڳÉ|�h�DDZ\Ũ��c�/�H���A݈��D`��-c��R)X^n�S�H{��q��s�)%�\�u4Q��.������e1� Mc?�~�)��'�3��BϘ'��ڻ���d"�C�D�X�2b=�3&��J!�ld��K+���v#��[ ��c���	�4�q�a�����o���F�/Y�\!ɾ��EǑ���c�Ƣ�%M�A����eJv�M%ؕAک��������2�v�9����?K�Q�ܸ��b��^я- ���V� ~�~�	�f���]��{pay�����}����r�t|�`�;���_Ɖ�}��t_N�T("u�a��$v���NU,�{�FS[�������e�U��X�Wf��ʨѮz� D~�|�N�澢��Ó�����U��P-��X�1�/_f2wy��ձ^��}��@����7�IQB�M�K2J����W+�eE<TP���@��P�� �|-4������HȜj/���	jt�;f�é�h�Eױ9����t0���Ng.��d�Ɍ���#=���1`8Y:� '��b^�SAv�=av��b;
�|�}6C\��(R��/\ˢ�c���1=#ZP8���`C�1��e�A[�ϛ,����0����4��sJ��3$�����R1��$��߿B$5	�͂�`ɜ���8-Z浵��ja�'����4ƒ/8n\�z��T������v��o�5��������ɔ�	:g�C�O�R�r	k����Ъ�2%�گ��u�4�hj�����AW��J��`��i,����<�@��C
�D �Ap�RO&�*Uw2"a(A�/������i�f	X;�W��R��"���Ĥ��������Wժ�~��q���y0�O5m�Y%#f���0�ڿ�Iso�w����hZΛ(0H��LQ5�h�:��r)��r�B�F�$�B��#W������l �ds�ՒN���Rt���7���1$'�Q�nY�6���YT���H��TP8�x��OI��B��?�}���:m���ܪ�b���2��\
�=�#X�H��=B/��V�2{����Ѻ3�:lvA��ߏ�����х�慬���ǁ�H�I���W�+0��I�=�Sa��R}�Ē��@B �7����Ƕ�\��w?�7�Lg�	Md��;�hS9�'���xW |�����+��%�I��Ѓb��WN	*�M ��AGq�[(V�����zr��u: ���0!N��Rc�c�_}b/��Gw������+����`�^X8ϔ��4�������4�rx>�F�O�F�K u���k��$�i��>�����"}�� ���}���`�3���|6�u.�|]	|�@_
a�-|�7M3��������q�RX�~��?��8�*���>!���>�"<�د C����B[�c�%n�Ut����. t��7�[K���g��K�?��+����mF�1²w�`+�2�P��e^2ǘX?�B�H�#Q�ey@{�C��^��KS# )�C��fgu;�/�|V��dPK~��#6(&��s���L�3MH�
��V�*�j��9�Lm򰯮����g�9?UAo��g#^v�	�
�t�@���-[@�P,H�ڬ�{עth��۽����|���t-��̾'ڿ@���%�d2��+�?���<�W�Pk�1�k�`�ș��m��/0���u��?Ow>HD��i�غ.�h0�&fy�5^�ﰇ����,�^!�hD�n�	��sl��*u��1J�F��e4�.4-�^�|�C��c�������AA%Y��v�bR�w��#+󖠵|��59��b���>	��Kf!nxCF��6���{%'�L��t�6�g��Je�p��]��s�6Q'L6�(�D'�1nx�ġ�����q�$�W5b$���J1ܩ/c����Y8���dQ{�f�)�Q`C?z�_7æ}��UؒMs 9\��V���3~���Q���6(7gCZk�H��5l����M,A�?�6@|n�NG�ֲ�m�ׁ�f��I�G�+���O=�5ॏd'G];�J�r</�i$T0���:�#�D,KI��$�܌�ҐP3�?�VI !����L;�$`� �U�?�3GZW��5]�~��fuB���A�����R��E7T��SM.#� b���!gҪ�Ƅ�QY�"������j	�@��Ӹ�˳�1/�h�[�(t6H������.��n*@�F<�[~�U2�~A=Y��ƲIs�u|(���{����P��`��طTN�eX�����c �!�����ãi���]���N�2ӥ$�c�s��YD�a6�h�F�;s��<�9����JCXl��Eav��so$:��_dd��뿀j�О��0m���Aoǐ]
�-"�|>����.w �<�R��jmM��a�7i_�o���0�d3�̈́co@�}d�2�k쌨M
�r(1I���K�_r|�r4��tqVC�9�
Av�{W��e�$W0"���J
ɜ@��S#}d�����A�Y�c�k�k�²M�*u�8�@-��A����*��36/��!*��>�q��N�����0u���h�Q%��|<�t���k�j3��)���R�^aʬ�T����l�-l�,�e^�yҒ��+Cdk��4k0�UjV1e������޶�}�ݦ�UyY��8f�|�dB#��n�7���.q��C�J�A`VMC�nzGՂl�cYx��L�����y:/�"�n?X���r�#d���ȸ[�Ӏ�*�܀��x����0q�)i����y��x������!o��.7���ʪ��,�ǟ��ҎS�FM����ʛ,q���V��F#l>L_�50J�X*��/l�Xw�,(�����
tl�E�H�	1^ǯ��?��P����i~(d������|lCw�tW�f�4�u7�
���M
�S$qs�JR�����׀�kFD��Ԓ�7�l�]�;���/PC�U�Aa���I<��l���6r��6�5�$\J+M���>��e;�{�}���u%4���w��Y��a��O����r.��*�o�<,�o��C�c�	��E�>�}��z�ɸ��4��6d� �y�6��.Уbۥ������]:����޺��	���p�)�B�����KP!5�d}V��)�PM`U?��<#�J%u�y�
�Ʀ@R%��8OV�h�~
Ԕ�|~��H��%�o�� F�6M����%˽(�ı�s��8f��p4��.0�����8j�9;�!k�1<�ZI2�7\�r�B�0KS�ޙ����A�S����'\�<����B$���;~���J4�0˯r��^T�8OAȮv>��ṳ����e-z� �SL��E� 7�6��%{���q��Z(���|�#K����߫-6"�5>��^�bO�̚�H&NvTC�������F��@Z�ݺ� 2ƀ�`z�ܶ)��AT�{����o��oi�}�6�EB�R�j����9�9|?,ʀ��?�Y֬!�>e�'����+ �rh"z�6�w���Z��~ҽ������b7p��R��3�f�.�;9̳�����A?p}�C�=؂3��`�O�����B\{�fʕ���!�n�?`��6��N��Qz�C��%�O�RN
�%��}!�N�>�#�������7�8	�o:�gW�wN,�؜���X3!ߟ���+���'�E�T��Ҙ����m�=�]�E������wD�:�9��ƽ|�����A)�]Z���pD2��>^kmZ���:1�����%��C��P4��ސ��o K�GU�!E���뙗Ӱ/�� �];�!陇���� �\�)$R̮Ӽ��r@a�xa%'u����!L������r��w��i	����\�3�fc���4 �?�7�~Jv���	���P2���61�G� |��/9V�p����@�p�
��hu54r�R
� �;���R(��7�'{��w}<Q\��7a�I�ar�0���&b� �M<�02��t[q͎o�zatR��1Z;DUN�����<(��q38`��P��z�SC���l`o>b���(��1�Bn�E]:v�Ⱥ'�d�L?@'VZ�S�#��e���l�cM�Tﰭ*���"4s�`=u=G����RT�x�v���nv����t�x
�7��X	_Ҫ�����L>��A����O[Ɠ������o��15�0L��c�B�m�,�&"7��.��I �̸]��������e*�ow<��okYo	��i�Z�nY���$'h�}����a����ť}�s_���Aɦ�~	��lK��R��R�tF���]��@���n5g�V�m��T6P�I;�  �Hg� ����C�]WaXר{	����s�yOv)K�Z0�FU")MNv����	�jo��;?�S�<+��?kT<���;|�m\�F�c�T�7oR��T��]Ʒ�._��ϐ��:�B�Ob�1k�}�&0|
�an���Z%��+g/����k�x��xچц�~��fe�����S�I#�e\��@n��d�	I=	�`�[�L�{��u�ԓju�ޫ_�ؖ��\;��]�oѶ�_Pu/yf ���\N��_UFn������\؈�ŐO��nt::&2���h���!hTL�aWu:d��1���ԠME��qC~��8�*uM�[�e����衿)x�WD融�Z)A�ն��Z��Rl4e�ʨ�2ҩ���4�q<1I�]0�r�2�I�J�$:״:�ټńa<��Cg��y�*!�D㔝��6�.25��|$��5�p���CF`fN^�s�E�yƘ����W)xL�ݖ�aشVT����U�L��7^��l���&X���������m�=��(�E~�pH5�Ī���rv=��X($�5ˢ�Ň{��Uz�,#�g�E�8顇"����!ד�Tm�nY���Gx~z�Fh���s��b�q�P�+HNZ�w 6�'dk��䤮K&������������>�8�J(�z�r�Z������d�;ݽ�;�$,A��	�������q���8�K��]�#�j>��V�����뀩"�%�A�j�l�c����/Rm���� {�?��ϼjGWVB�,�8��B`r�?��T���L�n��5x���朘�*��4~�����a�a ��^�u����*�D�K �v���kHD��2�Ы��c�/��Ԏ��a`bF����I�.�֟�s� �	�,uD˽��n��wu��Ԯ��ك�AhQ�/ �L#M�Fi��L��HGt���
xpv�?O��Wڴ��0C��t�ۅ�e�?���4yl���hGFD���Rb)ue.���X)/;� �=)���>Ϥxw���|��1�����7�	�1�BS*��w0]�~II��@�a�Fʇ�rÿ9+���.��nHLn�V��(��[�~>!�z�[d$�܁2>�-g?=e��1GSJ$�rJ��[�P晇�P��{hM�ũX-��	��u�ia�lu���a�������x|���p��Ŕ�c�����ˇ~�Q;���R$�^)O��%�euT��	����2��u�I0�vM�:1-��CT���gd!��(��L�@�m���7\tFyC�Ix��_豒���i���=t�u�1��!���{�&��$�y#���F�	]cras�9+7J��z�f�Q]��Z�P�9����J?g������1����ۏ�i�";ɘYE;5Y!���˘l�c��G�"nxL�S"��np<������#g��뒻�fϣG���f���pI���M�����&�4���&��L��n?A�u��һX���Eȼ[��?�oP��VI��A�b��p)�U#�����H'��?
'n-
�9�Z�UXH���o{���+����N��DP,��f�����]�y����M����R�T�Z̭+N���q�QjB��.��B�}�����L���:�mA^�4ܢf	E�zco��{�`��=���4U�[��E�t���ݙ��nt�M�[f��ʐ�g��I���f3׽X�fk]d�x�Đ�#�m<�����I���I���TX���G���І]��g>f�"^�k�CY��� Hcڿ}�&�ߩ�v�����D��[��輑u7��DP��>�?9ؘf�p���G�K�QDfM^՞�G�?�ͳ�(nV�\��D5�oy1��s�G(����uc�O!95��aۉ؞�>�je�3 4_ˊ�������2R�a3p[X�ͧ�o23`a)�\jJM#�:G�����zP<9m
;t�߄�P���އ7�`��h3N_2E�2�-e}/�M_�R+����	N���InnB���jތ6�#k�:�� ^]����"6vh
r� �}��l3DN�Q֎����h� 2�G�0�=���[��t�#��<�o��W��!�ĉ�J���y7f�5��	(q�Xs��#�� �V��[�4��-��{��HX��ѝqx����j��ii�4Tl1h��rL���*�J|oB����Jqb��c��h�7�$�CvQ�tl%�"hlHq�S�H2���zf��S���/���U�Kr���sE����q�mT��x�K����?f�k������s�Hn�-�����B�q�:��h)�r"�J
<����y�7�^������iú%�٪�;�����Ƿ�5l�S����u�D����&���(]}$�5��.w�6������)o�n�[�v$��;���(^j�����H�	#��(*58��)K�����,]�1��!��<���䂇����K���Z�2�>�j0ڰ���Գ�j�ai�b,�5�1|�!ttj�3��G�s㩍�m[�kJ�W$���O�`�Vɣ�Ď�`�eLt`���n0�*��%�Z�4��.�8[��|����F)����9�����b�Y�T�ͧ#^��<+4|�p��ﲧ�^�3q-�if-��V��������^m'�sؒREU4��շ������)8��c�e���J�l��|�1��,�=v��K�f5�W5����(�W��(c��F��1Ȋ�$f#[��|�*IF��ݮ��c���Q-�!+��߻�(fM�k�}Z�Aq�������koHa��2�J0t���'JN���Z�k�x�M��S4� ��b�;���
J(�N���5z��lj���lpQ����̗��BC`_����W��0�R��v�9�/k���y���]���K�O�-�i����,���Ԉ'_����$?���̪�t4����R�l�����T��Ad�=�"����;��Cg,ѷ��.�?�f��Pv��O�vGJ�ECn-r�uS��t`�����ސ
A���Dh��*5�[��֎�2� AO$�Re�����/�0ijZ�Jsin����o�D�n����-�|>� {'�)��f��:O�#]�R���>n�� k����f���i�nxc"Q��/�*�uƊ��܊����Ȣ�70��F0&��l�@�P�Z8jv�]��iؑ E���DȢD��'��Ûo�.��u���o-�~0�e�Ɉ]��ڝ���;�=e�{�� �}�?'�@LeƎ(d~y���tab�w�:VG��DE�A���ā� �!9U�+�9H;\��pз�� �`=<�Ҽ)��B#r�G�a�V�c0��Jk�ZC�����}���Ҷ�,@��l�e�a\�3}�z�샓�����"[�-Dh@�ԭ��*a	)����F`���a�m�~��c�`�ә+ N�Y��ҩ������(q���T��k2m��X����&���v3$ 2�۰����x2���|��`�e]���v\���Ꮓ�Z1H���ݺ�q��<v����u��T�]�W��	�)Q�=�t_�+F�!��Q-��,-���+��
9q��%�5�r����� J�B�Q�ֻI�����n��h�kA�jA��y>��i�� ��}}�}+��H�oxQt���6_���^̜���s<�B�����Y�HtX{��m���� k�*��:�V�MÉk%�a��I<�&@"�{����ا��ҩ��DRMۄHQ��T�/�zvB�4��v��������L�@瀖a~��R�@@&X��8�6ޤ���8���A���3;�
 +���Ct� �M+|���	�Z�(������v�e�O�IF�u��N4U��N��njw�C@4|��К�z�gRjWS%�y�]���J���wa2����0<+*T��#Ao>ѫE��e���ER��� O7��D����2���RL�<��d�X��o�?<��چ��������:��#�Ȟ= ���dD���>Fj�O1hei�⋕��@�rRr�/�]��J�� ޖ���0��"�*sE��-�j�"�+���)�Y~̅�W�A�^�����خ��qd���;SL(�$�������J��yxWO�%�3�<$ț�)�3�tN�ӎ�>��.K�NZ.QD�d�m����������
��\x�U�G;+��T^�cc��K������4h�m�t�3�� ���ƀv$�n��_����ϰ/����q{�H�s�Ũ��ŰG[XV�fO��Ev�|�iGY�B��l����fǒ��T�xt��Z��M�u����mߎ�M&�7TP�gN8$E��=�v���~KP�4Ps7
���s�*ƶY�����ǝ0�W��0�x��4�Y�)fT<a��Zts�\?��&f�5�G�T����S��,~
�m��{�h*iP��=�
�|��5��5���=��q�G��_�˝�=�&��h	l�P��gJ]NrKqa��+���L�QP�^C�r�Q�AL7"����Q6K���~ʼ
Y=�,�M����F`�_l�l}<S�o�����3=hXy'ɝ�P�Zg��~��hMΠߘ��3T�g-��VS��,�#`�8�<'�`Z,���[P��a����7���]2�	}*]�cxP7�Mf���z�\f8���6֢ �&b�#�!�i����Q���cC��M�3���uvF�z�<kr�D�Tr���TQ�I�Ғ�-�&#�fd�k�PMp��18���(&���*N�
�J"��k>�  )E�F��{u�v��r4ҦE�Ѷ���
��7W�*�$�Y��Tf3&\���� =ܱŀ�jWM�M�))"�Y�W�[X��6\��ҩp�k*^���/�������K���p�ڇ�,E^$ή}�!_�Jh,���K޶WGvx - m��Ѓ ����2��ll
r�������^�.�v�l�$����c��k�>]��E��Jw/F���Ch�۵���;��Q-'z,�+z��x|~�Q�%�ж�Ñ�]d��]��$��,�%��Ѵ(� 4J�zmm�
[ob�[�l�N���4	����_|6ڔ���1f7KF�FgM��ڽ�:����*��=y̐z�^n����5��:O��}�mZ��ܰ��I)_��L��]��.�`��/[(҉��񎱝�˪9\r�.�m_D��t=��p~��?6��}����gy3qs��)��cx��,����s�a��|��{0� ���B���j�
u�ߣ��^�-h"H��m~�}��'-ܹ����e!��=���U�,����r*Z�E���P��P�a��sbS\��|NMc�z���Ɠ�w� r�&m��m�x�����N á�i#��4��m?t������+���z٤�����sEx�0Fݜ��Xt��g��g�1^�P�1��*P~j'��k`X&L�h�|Ԥ8�|�������C�V�/O0c8�p������|ob����H��'9Y���������A�Gj���M�O@�����P�����@~g�������S�ED�=�mD���<���\�poq�;v��:��Ƶ�G��.�ӈ��ԃ�-zk��K�M�?�k��°S�c�v�e��m��K���^��,G��L�:����X��K-���Q�>P����(U�*D,@�2��2m����
�<ٟ����`
��s^9{���
5��귵�|�E�h{� 1��G���%t���v�"_aYŸ���N������s�aeú���Țz��tWG%��@D�� ���d�	�߼q���%'�OhCp�9����%�����R�Z �@��_.�]�|Ϫ�OT{�k���$��~�����u�C��?�)�/��8�*����}�M�[ܞ�ȡ�����\e����0��𸓬Y�-���I^�%�1:�f35���z��v�  W��`��n�A�Y�C���&�f"Z\Y($��`_X�"�1ڊXP���m5zr�/nV<0-&_��xP�?���+}�}Y�-�{���Y&�x����X�Sa}{���(�J_�󕲸ӧ])x)��d��vo�	��p<��Kn�fܩ���AatU�z\�߅B�49�