-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
N4gghaRTrPOhVPiKksQ4813zeq+WAUaeA0bBdbRRse+nxYPot1bgDf0KkI7OJS70zf2JqSJF6Zjr
YJB+VjgpRpXxgVNjPSqmWiUriw8uiOuBEN4N8Jus15v5WWjpgBq/1CVFzBiZPETzjjs/UK+be7KF
Nc8Luu4X6ugnTEs03z8X/HSFGtY7lhBSgFl+08gupJ5AuTSb4rHvzG6f5vj4sj4/t1qymtDr2MVd
bdptMNt5IE1iLUQO5fVdh4ezyEDePmn6mtYE0ko69yS38igKVGnffgknnY3qna7W/1UMnHv4hngz
w5gx4e5fISBHPlyydGeTe9dm37SC1B6fQBH17g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 49536)
`protect data_block
WNBgVyZkZRVrzOu8+10fHTo7wt9YPHEN1WDQqTI0w9JANRLmhCFk5g7ItDi/teivT6MaHiA3LUaz
DZ713AHabk0CRkDNrUmm+7sSSrNRq9t8f3b+3bPgMR7WNBi6kmoQQQOBG0h7v8RnCggcGaJR1ais
qCPWzNjgBi/oHpmA1y6tH/q+mjq/FoQF2LOjR14/6nwPeGlOzyBuDvdsbKZ2hlMSqxhoVL2D2431
sHLRJea2xGSgd6Ggjpl7S0rzqGQKPGgUdXn6JGhMnwopjcRTsEdWbnQz3WIWkqZWfTZCbCrZ1c8n
cEJucBAqZkBdnTmIG+Xuj8VaWkiBDE/k+CIrKrjxMr0sSdBRkraS6LM3GaAub12u/fdDnvrtohOw
Kniq8Hc9a2wDm9arZ6z5yq44ceUC96AhBcARfi65GvQVckxBvqk6QK3/pKSF2jRk0/vQ5X2W28v6
wOWjG+379kxd5Qz8LSDee+hM2zxmL78NGKic/yTPYsCDW+y0o3kxdLFwvCp4XZK6oME3/MaLzI8d
JouLg/gOeqwPfrsyyWsoI67h9nbyz4tPm4GhLYYkQyF4vht50cryZnyCznI44Py2lmlx/Ua5BZwe
nbELTsUBw4bpDwj7/BVZ/XXdDND6L6D/Scw9ElEgivwv0YF+mGHZo0F/SYCzBPOhZTIuWOtZInby
f7VXRI1qc6fs1pDbmEk7lc/7w8SVCKYU++Y2+c+fvHfPN6Oxg9hBdbqoMrvo+DHdNRfTCdO8Rq5G
2K2XgTJgKUeVr+qhSwXuSuK6KqkAGHWMHYW5hqjmm9mcfV1WYcZm0/Nv2bDKWT1RVNokOeFrOiAA
91SEnizj3y00+dUrKVqzAoGhpvmhsb6WsQWvnDikBmtpgm5nkEibpXfel0IZfD7dr3XVWXIw2MEp
CwoQAFspOtQtrvvSqLJZJ7k8YjMykIXfZsBe4fwrbAvqS6DhtlYeqqofktkyBFoQ/ayvjG+ZNPth
JyUhpDsbUaP5ko2kRQEpuQ42nu+MOVbgAUc3J1MWb3lBAY8q298PqZTdFct0+eNXGQjYJpDmHDUk
2au9lXg+OeSxC3x1Qp+S+KYEHl2tcg57h+Nexp2xbw0geZXpUYi+16WzSJsRlLPa/DvTTjB5+TCN
csYySrbe8HQJGDqGkv1m3xovvdyb51erXaMP2lKCk21YYdpnek5OjaIl9eU3GVtMHO1SB4ca/dZC
dGdHIeHd6qkFRhN6Ingj/YChCL5qOapS+eKlkTNH2FyCiOPsmC2Ly4dGRdweuPDdMcVbg8pS/AQA
YvFU5czIzSoKFMtbR2lKU5XNpA+oBF60z1oedwy0wxcjyj/p7fnOKXRJGF8tNKABCsbvgBzUReLS
dD+5S5onrl622sxgPxomWhuvZvSL5X8TJ+q3V3LClvEmOYnUA7iu6usedQMPUt9y+OVKRq+NHb2+
4Edrwrwk6tW0vGtMeVInpn/gJrMZoOQdqmuK3XXr/7aROPRFWGasUU3aYu3RMnuscQ/gJhk4xX5h
8BCwzuEXedufgw/fWMW+LtsoEqQtBk93VRbzV919cIqRmwDzkQLDmRg9HDyRgS89XhMOEjRxFVZL
rb1Te9kFggL6mREu2DA9QJRgiq6ArlEwVhCzDx61zNWIXcrOdybNQo6njPDC1D64JI7IuG5uiUiE
gjrbopiNyQEb2WRHTAPtLDypDo4RW/D9Del7mur1S9sZ8Uh4f5CtsZk8IHaBsuA9T3CXC+jKoZWO
aJvG/mtWgteFsw+0WE+RZh85IWs0yikFNYVW4TJ1QtxUeUWSLjC2KemQBMsFJ10BStI+kL0994E+
WoDDNWTEgR6Iw+cOew7fKIIR0u1DVE7IFvgvcCr7j0l4rI90nTdCi0Yf4Q/ayS+/HXxrIRBaTp8e
jBtjO7WbMk3PyfZYkHAm1IGTKbqn9HOqdHdixBYb7hF7u2lpd0SZ6Snr+HhIGKlL1bdsw1RttqNu
eRYRuXqvAR2teqzdMQzTT57Y5ylfaW58/BMcRmjs35sh1YPseAlFoVOiRln0SMjD4o8s53XQaZcg
46iy1VWlLSupD6sGByxS+ObvfW44nWnZiBRQfOnFfcOSPQSRkGY4YTm7ndxCq6apB3zGT6V0STAa
zP65J3yV+QGX08AJxRY/DSnkLx8Fo/NCoXjk9pIhdi/1Z3RqQQUe8sQg1PrsNEMfVRDKOpQx4wH/
zX/bMEfk88cdIlZOcE12n3yeRsV6gZxQd0etuKaaTRjdqB876AZHxQRB7tIKH+3Psqv4ibHo1SS6
CsrpQ4ckxhn7c0PVBP0muwFC1F1UG2Tvrlnaxrqw08uc4TVC0uEuWfbYL1XdjdwbsowZRn5rQNED
LsbW265jKEFp+aIPE41pkFNBbcnrmQDrJ5yBNPVNygI/pF/MGMoTDmo+fNz2QjFL96MoWkyZG+xO
hxqC2tADe0ACwCyXVZulZAVN8aKYX3LZ3PtIXtaeMFRcAZdlnz5RfnwVK/o28v+fjkTZd72iNyoY
WkBGGmaehiZDlt7ch1Tkx27gQWWE65b66/ABYL0foOUO6Y7+7HKrKP6kxOrDNHQEQKaVff9tAWLc
5NCWMGCmCR8gekXnfomvcM1XVihi7L0zsuKvm945nDTHBWGLQdtYPChAcU+C0zCoY+C+VemEHlx8
TeyjKJuonWXYEedxTNV+jkLLRf9EBpPWwT2gbtkdpwn/essXA28x8dnO04PtZxbQlXWD5wTmpoI1
/GFgVZ1w/dm2DiRpqLud6o33fG8Qe/t1RhqOh6WhAMoXF4hWoas+CuKbi7WMPlYjaARCoMpD99Gs
v+tJQGODFg6XrlAIRNHCHcAmCHwVFHrFppTa9a2pYVl6Z3y/5rKRrgZasN/b9Q+8rNp88bQUveW/
AiEqPeIJZcePCaNehp+UOmwfjgx20aeq3wY8DF+yd/She4t9FBUxMWLHI4D+jw3upeFu1SKXmav8
CKTxFBnLfBTUdSz2m5rrRNTOCHXKGX9YPlyXLmFeTC+NzX+Vjlc68khzsrCfzQzExrHGLaFBAYE9
KvTdLAQhEsou5JBjXIHj3ZY5E/MJmy9cyT6DDXU6DsZixdPiMM64JUGW7Jfjv6haBslElv3GeuWn
d/RAezZiLCKKYnCJ3AxEYLD7D8nKA6BETmt911/6BW+ROl9GX5EfF6wyvRDcpNlxgd37iKUmomIg
mrN1MePwkuhHOh57CI2LrNsHWj7ej0NWssqAvmOBX7Ce0CMymD6hpn3fM/0B3nY6zDyvcV35Z3Yn
mJon5tyHXoLEkuCsybntZFp+kOzml+ELkaxALxeDIX1IdwujuCb2R25EI8TNIQDC+9o4anRJzY/B
v1jss6f5O/yZPRyWa584p3+HAcnnY+YrKkRuRcJ3FsRCIgnKGrUL+FJSLkNA4w94Sh9qu54+9gnD
PQc5ea3y46X6rE7VC1wlJ2Wikts52XBTw6LEBAo/ukeO236uOyAlPwnnDQDz7OVHXv0Kug+D/5Po
0QuKKUVnu85RgQu6HjOyNKVM23heOMfkFVSzr3yMXLt7o4+w3UY2CA+8EI5twZgFIi8xUWHhhtUB
WMU5ds3i6othH4K8UKBJqK/7Ug7QeKxvBSduC6LzCIXwsTNLRtIc2+Oiis9QjIbhawaMR8lIez3d
jUnl5TWBaAsyK6VH0GQH6k/Q5AgbW+5uYYowa7NytJnPn0XVUdWURsLFCLW3awreM6nrnNXWNp/R
aJ6CqeanQLkdFK1GnYZV3lS3rosyslfo1Bim+0fIftcRPL1WEB3SXaAL+85Ff8oPnG/UeCq7MdWJ
sQpl46iw6jxsM0m5dGa750I/qu0utC5ShLnd93VUy3XGt1tkCauFT7bJDT0B+YsKPXIK/PETHJhb
kGXfMpR1cIwnOcYVcU3DAO7p2b5G4Rl9jkDf/MLvfOVjS0ih3V+NjAR7iSHOdj0yn9YUH2IQUabY
I/8yFM+0kANBkXF/p98UMJUBfguP0UQvHn9CH2o7BvtIx6FGoJ3iUg7ae6F7TixfzSIt3/9T+GTW
QIoS36OmUmoZfLZCmN2INJ0vTrtfijDYIwbGXamvZodMRkvEsWojdpko/BIyRdvubQCqU9MAsmoL
YMO8IYGF07KfGR7y56Eo+MQ2/et9G/XHbfWNVvwGMhPI6N4CGisHW8RrJcv3zIiAW7KGEkvwftoa
k+01k6NogmJxfdf0afOryZbSaoNsK/clWKYmON8UXppLsxtqU/ev42DniTFN/d0X0gtoQ+L35TK5
xe8rtwuWsbnrTZ0Q/v4N2gaZXENebFXAUo9XAgGUokr9wtCfGtB81N8s53tN6IGTwomaHh4UyXKM
UV1DIWv0HOp6kZtFhcuRa5TOLwMgFRxCIbKF+FYpruqqlz3yyWSpoBIfZio2sPQZP2XZupAHojtX
sABRlKiBamml4NMMm0A69efZ2HXLjGoGK94zDJyMLf+o7v8BKE7HaniarMSLlX1VnKeaNwNG3riO
B1/j+zG+KpdnRHEx4rsumfFZDdyev3G80uCi+DB2EQgnsbvwZN3YyyvEpoLMe3/zcX52Bukzrggh
zVa1i/tp6WNxdglOnDFbqFpG7Ju/zcSvxAaZs7dYoVjbL3y62wXiHS1aoi9NHj2Golg0alPP4ePo
iWQt7JwRJPQVZ4KaCnblCkkgidNYGP+W+6oc6RPfiDyG0LKkUve9VuEKbley4njTVXFbXcIAl/Rx
304Izy3Lu4hBayPb0kgTIbGNOeKU6lkBDmNmV8sQhwTjtKnnTCujGajsuUdb9T4GU7Ssp1diLgdn
uZNt+xVJLX3nXIkItei7b0IVurdckjXxnIyFmqr3NiDqxmeFc/8Bn6vkTSNkyF9o7OW8WtrHDg2e
BP0wELyoxi+t+tvi/eZrDFWBj/G/vmgGmCPGEK17XBkSK856H1Q9d8Wk96hJIVMQoCB8xygsVOUJ
UcFwbQUOK+3Y95/Ma2rYKa0Czl3agwF4vGxvJ1rIaETcc5RBwUpeeE4B5t+OVBnwHXOOyrUz30LG
ck5u/J1IxpR9VWrDziijLx2yA6lKOg9zh2Sc2uVK5IC6xYgdso8wFuGrJNQNdj+/8ETogdslgwU6
Fv/XoqVeBCZX+64vF4dt1wbmjJq+VAjAfAlA99QxIKs9tWwVp4VOEdm22W3T4zrggYGWKoPAKCnk
jLXoVfWGOmg/cwMWm2FBgVrQRLbEhFG4roc7fJJN2PU0dXylLSrKdlCbCEDhJAVPF4/gjCJzoF9q
ywwnJgPZ5UVnYUjI07D8pNzEJ1NccXrlBfeed6bJy+6B1t1ptsbAYN2R7BS/niaUNqZcXiozKZyI
KszuMQjVWhmAkFs0KuEkIS3cguDPBsWITNqIyjhUebI6DELjUEwQeqDIYV81uAY3KOL4SvNNNnQu
e5mTovQ98dpd8gUUJ3kboB+ppUKLddY4UfhKp18xfWLbUNOz9UiZhZpwcjcO8gNO1mpGLFK2KuYy
Fcd1xW8kf7+Jr9d1/3oLIXWt3q68USTb8zTTC/srf6Kkt5kEQL+g0LQz4tyofgP1IJ+s+t4YVYhb
LqMxzCGGwLx1sSRPjb/zSFUOmbbvxpR54aI2grcSBvKPxhvVI2D3GOjebjrOJneJwARrfXiyFv0t
V63k6L4DKeH67pWGEWmx0gxrPbVjiLJ1TAFJM944/hJKIjHUDDRCP+LFTpx9Lbo809/Ea9J6JExX
+eSeT3lF5xv3Qzu3B4bnrTUnHUEM7P+AUheFPlnR4+tXjhMGjiHwb7e7wXKyuywI84s44uiv9fRl
KsICjrts6iaSQA/9znpJE0rMrktKnUwn8K0ugtbZTrQrOkFfoA8Ps+7lW36fpkbqIVSKBQNBj5wu
spgz9GC6nwzd5lN+R9oNtY/5sF9psxMzxRBwUgU0ReUYjFqvsfrII1UIDWGytGCtcVdXfSRT6Z80
/fprGXZ1pBk7Tcc76v9fiCTGydBiD7MFIf2R/trMZMYvpK6X0kpwuzrosdM6U2sB3uEofeCNPXWp
e5WLkbxMlwMq5iw3eXGvbCkpdi0gxFsBrpptsNk52CD/1V0EXLjDdNF8iNYb7HGX0k2cLHSb6oJx
HEsPrAYPwLvktZqw8hE5ghCqeZINTzjmoPeybTiBeqJ5D8hp5jug4Ydddedxc+TB/Op6wk4RKJOO
ozoMUPSBwqj4Eaw/nvgusjVowNxF+ADQuWnjpHmktOY90HL5w2tLdnOZCTZf4vbkb4jHltOPyFZg
tNu+P6vIK5/TQikwyKTlF4cV31SxAZMq35wwMikWCRwgvpT7KrjvePEP4AV7rPA456sJ+DTuJIZS
nJww7oCUHON/deRqVebWjkkIkVXOW4xeIv+RrLVRMTfdok+KrKdnDI854jPeCrtMzcC1reZ/YJnY
gxRiFjMeVLxRq+VJT/kdJ53sYnm+A5I19aa9D3MNrVXzrEje8RXRdEPEGoEfh8Cc6vol5r8oX5IQ
FetfQI9+E3WZ/rxHVOLlgVs0ZAkSJKjtMGxNYzuXAb0emiaGZ1FxZVZVKL6P21vHZ8NtkaavJmK1
Lo6zT2HGHT9s+vjchudbr1HVjqNsLTF8cP/P0rU0cEQKo4xs+Rk6y5gP+OtpwfPBDWFgSjw7CqGY
dmy3k76/8eyZHRz2MoNY1swlwGdIGhh8xbO/yhXJHUXaZbFc93JbW1ywSHGqnak0us5LXES0P6KF
tn/1Xn8CGhac3T6o8Wv6OlP+Fu4kupcttuqWxMlQs9IEVhvIB0t/AeEOcSByxdaCR6L9zoRAl8TA
6Lzu6D3IfR/9qdN5DgVJq75jvcxHHJ/yZimkZ4Doz+fPVDNd8PiLKZ8Tk5qrqzor7uGznrFIdmKn
netJ1bE3arn2iu8Sp8t0bAqQlYvG1E/i8fvFUmNawdgd9HOTnuasFsC2i9D2Xyxr+hZplHeUYjTU
HzLqPVG2L04cx9EFWbn0iL7KnfzXhONe9BxOT9EBVgHgRymqmAthvDLHsk202i2jxj0EF9R7RDXI
9ccnUugHY17bF5L1fa4jU7B1AGLhjZ3+fKnuMSY+3L0VeUeZAZZhACj0aCB/LXYghFtoe8VOZfDo
X97rxgCHckM2Jvzc6YAURiuiLf6lxxn3ZjKF3sfcHrbsYdwa0ZpD/YTZ5r68e7zfqoQe1hEguZet
yBT+Ia27ESnLiFj69xz9TfrLyPkFGx+YD58sqK2+iakz1F55e/pDFCg8ZKmHxQ18WeYWaK/rfT6k
sH5iczsqWFiGQg2dw6D/zeS2s9KzDiwGzoF2IoAu2cbcYjP6+EU69QjVuuh0SveoAqs+Lk3udyvM
erTc8qzGawUDNvn79+lyCr+n+RhD9R6hmzB2U/8fBgqK3d3oYs0bfo3BeX+SiqdjpMVIuBnuYGsR
uh/QsAcebBexdf6mCjdTAL5uUHKGOQvQsQRuVBjZp3LSXzcsk+he+2KIxpAbmID75C11lMghK5dT
1ivUwBPSGgHDLOdKL05eeIbcfRUnvJWGZUXnFKPWuLz4Xyzx52n6IrUDKBsCrrOA5+uSDEf54qiE
b7SucKRba4TDhiX+Byvdg5TtA9NSIIvxbU73G8TzfcCuFh95l1QAcwzISKK87JVbNdZA5bInhXNq
znhbUuL5pb6VGbakkSSFZK1CUh2rYgOsiOEl7TUPmd5AZRjjiAMMyrvdO2jc0HvPImdydSLZEP60
0MTzEN5U7LyRdGG6ieyw9jwR4SjZ7Yjzvm0SW3nfdfbkJJ23OJovIpl+K1JHBxXNL2fUnRWbQNRY
7qk3abEuDjAzSqRq/gMUVRojUb5SfO01/jA5+3dqaHdKTVE6N0ZxsU9vYERurjkiRmGkvsHkSFCB
5x6HWSY+0lsLT+yIkKzpc/J32j+lnzL/JVVP8cUQl2Cx+2AwgUjoN5qc0HzxpKQLQK6fu1i8j/Fl
Zpq2qAc7YtBMLj6uu5Mubtni/FGicKA2++FDg807cIV5hjs9Tugej5JvuMFJQ4fnPEFXawuaksmO
C+RkAhQt4govIYekZ9QUeuOPHPfH8GUKAxMiBPvtHAxqiOiQtitQWnUGUQuyJxlp80YtQvsvRnxt
qTvRc9B6N3ColYluon4imhP7PlKKzDUs/0ANcHoVIKcdUyq3aPol6TOmaJ8FvTpQH/5LkWSA1Omf
9xOPAsoNqdW9vWoIZYkqnpy4h72sot2+dxR0z415ME3ONCebZuLmDaR4FpZGF+onNcytT8YGdVaC
L5C15SZHGqnSNo8TvCn1bseDk4Skf9pB3iN9zPtpqoyXMatAth2txTaLK6w8hAPZWBl/cdIiksGE
YYLJ95Ag20rggc0gOd0lQt3jLIRj9z0YhNHi6X1gRwG/sXFeAwk4vMlhP7XGjxxGqgIr2sX6l85W
L6AvYwdWgeck1GAgyfQoaPRu96KIwe8N6XX7W0m0PxVbEyMFGhOo6Tq+HAIgTi6Big5Kk0GslmXH
Vo87v8gjNk/PXsBy/Oa5GvPfuxNVoyA3tf10vPGOMoh3MeXgcAoRdWZBMNxNLbd/DkotaHOVnlqx
t3sumE0SL5+QcZhnv0zzPLscouhmp1c0r1lnztvNL2tSEsZBbToRgI+QmxNdPTgW1jCK7mHrAg2j
gLYrmpaVey6n4ETHFP89VSYP/TU6WrhTe9gwrGMxRreMkoNgOnFMJD7oo7mtpDkN9vYOX1Lz62CO
aoSbwlnTVJYCwifX/kkzM+mpsXy6LWCGtAZm9TScsbqz2bEOEW+uTgkOlINT6YYusCxkvCcDVsNH
9vE7xWHQzOCYdL4Hl17N1Ecy7FlMDAz62mqsrmC6hX3nn6CgVX/kUnrXPseDFUNRt+mSwZ0qaCni
MkmjxYlSOZVK+3fhyQv5FUnnN0AH52zJg3li1Cm1fi5Z1ySGaM3PaXfH5QzZFlA0XvnAuSOhc0mo
a9hSQe5fTNL6jbJAklnNGdrqs5mUDrUUp1qiyF8cu73BPp2SkJEwekSUQ/Tu9sG+avSFdZeS06QN
DIgYgKn5hmug56JrBay95gSfLkcbD1uHwQ7ZCgtIKhuxhuVEseaHCWlhm9I8CWquSGF0rR4i9NYd
sXOjT1r47gxeyUZzQVQwqoHuxM3RosZimx4kPpkRCK4m8iCUTaijyJJXu1uPWq9pDcjUmtfH8vbX
XMVQDpQ7jjvyeuzvqb3EyZ44zfvFoZIwwk0Nci+t5EqUAinx9Wz0CVWxBULowHtUntLmtKRo6RZG
GLQeMHcvi5nPypOuU0s+h3cArg1zxY61vcOhgWq+ylSBxaTNJu++vb2vWA16PwCbSOoVM1CwOYnN
FPGHzwzxOnMULJO50sW4WYBWTnVAGIoaGYy+7RqDwfAxkdvPSIZTOlovZsfNYEgYd0x6T+nSKH8f
cHOy3da3YUaxNFJ9MKXioNe1WVMIuzLk1ZA6ZhhurrVjR6I1anVoEOu+BAgEKn8C+NMbITn1nBd3
qgFnZ+6XH64eAMUwmftv4kqQj5Jsmf9A2k8mT7/resEMCgJAYvhpzpyn8w83NJY0o8a8WH+YB/Dg
wLRw0ytRv21Am5bWtPjyQ2NMF/x8LfcUGFH6g8ruQA3kphZPu8x32wcpCfLZ0IHHPb4kyqwzfdD7
USDLs6WZ9RvtQagf3OWw4EYU/ooCP9Pe0B2lpwpZtI8WYO1bmdmUrkxm/HjmsD3IlMCiFEWP8IcO
QjgWXCUcnvygKEXUrlYttMDI9SIlHH9jaIY8vl7F63laGv5H3TZcqnHaaOHn1vQ0u55l9UnLd1Ec
tR4IqEVcCq3Ng7ibfYAFA5X9WD4sn0S0HIvRwfT/vl8opDe3Zfc23U2Ck42Ub4VVN8HYeDJ8vj8b
xdzm7pXCgI+oDEOlwpb0IZyzNByQ8YiFC48T1zq5s2xr32Tranzsf0WQi1mY5lhr+GH0myTxXW2l
gNSRH/TNCsU1h7pvjGDvbv+QYg0vvoGlEs4EUoAIIq4FbgAT9pVLdf5ZWA5AdK4w7utdVYl8wU27
fDUoch0/6QKYLYZHgqMibMhY/8/3vC3bwTrgcVqHOXA71LXf+oDdLw0qBU7xpLyJJ2oveqaid+5U
pmVy3ifZLokVdbF/Ev9s/XoVALLBZ7INdtWfWHvf9N07AWIanwstunOiRfcPNlejyJ2fP60VW2GM
S5yGtRpBCDi/S9QdTlNfSgFTN3ot8fe044NrIe1khLrV60Qn7ynWAn6Cuf5WnWXzU33f1bysLG9w
WFrHmagygxaL+F9BWsJP0Zxy+Oyh3C2TEkSLCfu0msY/fxADgi9rcG4FQw0k8nzy07OupsB81rY8
4KN+1yfyWsaEDfEL16zq1jLNJEl5dY3ZmVtrIMiZrkD4SOoqMHZzJ1ekwCrNFf9DDPgx56BNHw6H
Quri9L7EWIZIQTXnwi2AoKk7FIP5V3/7PIEK00gHGYy6/GMLYxnoyJ1hpssmJCJExuIl/LRH7JQY
aTT+DMVzPrPkqUZiBWhsj7ZirveR7FBiFMSCl3RXPXVTi79B/P9gx4bwfR/oKKa5h48N8UsqS7Ne
5OG8SC33Wt1iASufo1DptBPu+7RclZNg+SrCSb0d3KLLSi3etqaYHbsTkAFe+9brsv9hjwHbDVj5
w37wMUS1CnUvPMJN3g/T6vIyC/eOqOJuhN970iqqh80ubfuWl49sCd9zbbfEEl/xxjWzJasqIYRt
t/Wq1yAiz8jvNUmJNeAN1oE3LWXap7iVVHActoeDNDHj7NjONRl6tmomrmrH+t+UWFohhmqDA+XN
/TEOzdK2ZxYd4l/CpVvhBa4fMmSNOGI5aeHzd1xGVoC5x3qXVjk1++8g+nahICmUKmIZxLp++ALf
d5DN3/XawjZaknzOsf0v2EpFdgyZya8kKqL/rhMwOhg4JQF3T4lQlzQa6lSuJQTXDldDiIo3Npe5
0r1lRJs7TLjLg1wBUGT+cAAlMyxb0nuzT6dQoMQHkVTBKu1F3Qnp5OWhSntQ7v/br4SAwn3wKPnT
vxPCuJEFXJlDXP9eCe28rSVqVuqEnc68ItfzVC8NlhSYT9FAAH1tL6fP7ZqOS2LG4XnMz3pwJnsy
MNP7Bmk/v8Jueq5khIEhYCpMQoNLOerhfsEdGuVeAsyYRidzkxu5IVFe250D6uOAaaZciiFArPmK
sTFcGmU0Vv73nIhQRN4S32NJ8u68ca4q1BVx7RJGWBkiMG42jHp2TomXUDlHZKorL/+jrTWCDmFs
9l2Y2E/SnSlu6M1Wyn6ke4LVaEZHvarXlA3NkYQG5grxiZ22sXFn2Cj1st3QD/+A3u2tAoisl8jz
KhpS5nXcjyVyc/WJVJthaI2O5cweMXxEMefIgf38oR94rzAsbHBqMZ3jpsVPivChRtsFbby6Z6pl
1B6rJknvlL5eaSnOtFeVf2BmChHfl5rX4PLDatoCT0Kl0hu72SgqWGq98NXf0oqVekC77a6Xdqv/
hITv+ZuiQNZf7UO40YpCK3kdC1Ax8F/AmBsyxe+9OPE1DyOnAipQvwxt/BgVmZKIkp92a3HaqSUS
WDRY+DrcMdUihQFuPlXYWSFmerUMSf4mY6mmn39D7DLVdsM3BNG8AUG+CKJWOmAPRvlkMq8EOENG
8ryXyBgviu6h9JAp632njgX5G8DfekmfwZyK5wTiCXL5HUhhftz+3U2y+/+04xRL0q5fQK0/aOcv
JChRcHbKWwjH8/3qJKy+SstLfxkLgJ9Tr2OVgffN4qiUK/q++0YaXVzn8cttjYNpMTzx78Q/yxOC
yfhjxkiBiNm0iZc0VG0lwKqlZkzkglq0ZrE65mqK4uTpsUpX/o5dYrr1hks1ZZV4vlaSSJvfLD2H
xXkT2nfrdBL1nVb1AqYQPb7lEvENQy+5XWSyF6sxL/s0nysH2Ba59YyUwJg3HKcqwBqb+3453Hoi
QvuMG+marBscaUQzkphRcnaZWZWJ4eeFyKk4eLTurKqTFEyhfmbftNhZXPia3emt6sP9jiay54GK
XT1a4RGwrZsee3Unswjs8DnihBWNwuDpRqZi+JbbrbV6YWjDjc2OioERhmvNG5+a2rEp8mQUBto/
d4WoRz9ZJq5toM2Ex+k7F5QqyT5o/E27gVwSi1YsgbkyDoKztm0WqE++tl0pH3ZoDgsbIAfbcY5B
8rqPmu/3QnRXIeCt62WeheAg19kJOVZwrwRl6HR+3AVOsQ9XvWnk9v7+n8GfhD7nFstMODNeBwCb
fPbeFamQyqsw4Xex5pmgxzoLs6L1AtzRcDKocx2BBPY2NDmDYU379IjHulhveP5rHNF2ARWTCg5E
kQU9CHReY3wPeOqfsF5cuf9K3D0EsL6SJcPz4oBIxdnJEr/boyhiJ73kt22qiXA4KLV+dogDF0uT
luujiA+/xQftaNEwM6GzlCdCQW2nSQtnzVq0Qds44TjQ8BhyC2Rit565g/eJXlS1s++Kw1W8NyDl
UItMiIXxRE6Va6ai7CH7JuXHGgy3vSQ+UP9bVJmxNbeqwjZ4A8EKE0uspIPfDt9g8iq+8ZanumlZ
3s+peqjuY9UxrYi0yK5N4gT9nUUwQW8wBnbErZaFocI1auoSmWxpRhX1WfTV6/gtxVDHe1O4WFwG
av2eMMQVWhCpVnazlqTR162lHRVjvZZ/Q6Njn8zzCToe0vaC9slBUG9RG2enbe/P9m7owOZGpuiP
XFYP0HGmST0sHSIxbsZq+9L5Buqq8lSCo5wwm5GEsH/RlZgvOCqESkJ1dz8WuYTm9GXLfghirEBe
qnBXSgv7c18rvQ6jQUxUU/XGkjaBi7wppUYv0xN737rBCWvilbvSmtmF/b94l/3Q0whHGyQurCOA
ZJlOKXyhTmZVURQ7vccTsiNg/tfScTFUnIbDO5xSAMfmQSquHTWDYbyZP5jljzUvx2axhGbzIDca
vNPdPrtrytZBJ/2CWPgaI0r+6WnPnWm4+Tex+w6AFHUHrYkRtHLf18xFJV7vCZiT4CE5QL1lDtdi
5w0TasGQHzq7gmnXKdPTI+8+eHingpYIa+pQFQwZNgCuJ1CcOg/1YYT+KDLmA/dkEV0JWN8kzZfa
T66WGtqPOs6zUbsWiSzCYsVkeLRizKmHjfn5JivA3MgRxALh2bT/zLeOrFiK6TtqOhvk/Kkst3xk
F5zsU5fPrbxG0/UbAKiwXBXVALUJPRNtmHjToF2Y/L1nsgTzZE1t7ovOX4p+lEbQHLILCPknfD5Y
79+BLMTRc1ZQY4CwYrKILer9681ULm1M0TTBmLP2M7ha3LxL1fDI3gLanBTEi4qQU9UC2otx4w44
zz6gZfl/1A5d54emH08Gt+ollL1QOpjZ4ONvlJOlhaLziBo3GbKieD7O4ZYCcpJIvE6uxhcfacWc
FdJDWjM8bTno+TeGuuHIyyx/FuTJE/O6X/KkeYs8lwnf2XEDIVslEnJzhF2rPQ/wKCjTEZwb71wm
n2ahK3+a7iWsZaqywhrNGhB+kVRg1u9vzoyzJUBwLQUlwtdKDbxwdGQ0kfzYm+6zCzpprsM+b3/4
QLIgh+KsVFWtW7Agx3BMfasqBx3X/gZqDjUM0kWDZ7Id8oRqXxsZOi/7NaWfpKEDJM9qYI0VcF//
6kvIZWb8ujLRfy2cbQlTkqvpiQG3Y2L/4ZVeoUZupeidE3PW+L2NM1JIoR3eBXlUdgmxfzIEvq8h
CeiFJpEJ297gfZAv3UV6Atx6PYA6IE66KDVblb89A/ngyUkGDTI962OkbWokZZirA6PeOPH8ONcx
uqE2jcOefQrrwsVRaAtvB/8JLV+qDTWUeH4xa0R+tRH9SMvijVeiH4r5ZrjyUeDC+M3n1YZEkavz
c8SXNvmTRIpDte43KQYBmIx7TaQUn5R/Fl5DkSa32dphvfZQ2ak54Ywb6Eq8LKqDNSZ41ZAcfz23
1dx6VGlYG09/CsWzCwbNINYdRx/T5eeMvs3vtP4Rq28JPNC2dG6412XnS+OvpB1/xJ/Pk50r+I3U
xCq9dOuSdbM1i2ysOUlSS/ETKu+zf0wmaYgSXNt1YoQZ/ilEVMckbuWtNBKJdtea7QWkYOevJBqN
+Iy8+iLxO0kxYoEwJ5Q9nKfZVEwIZpr1fWBPXDMlR3ID5d8dCmIy3JzKu2HZKLiWbHKs9NkAjAh0
kbsHm1wvx+Ho9SXVJY7PxhYZM2/ygjAeQVjBKR47WmR8Jp8CVOFbhAd/TFJ1VKFZNVYTmGp4glvS
zt11/3o8JF5t+bcDwni594DJSlqoI1+7GzmnXrWnDeEAT2BCw1EDUqmewmBeICGjNRrd10HmrHWu
A+DoKE57uKK9aJNu3EAih/xV8bw6EqzmhstVDDaqTr9c29abQUkHPJkoWE/8UQTTsUnovrkf1kZh
5yjOw/mOMORJZLg5BlbnOtTGHncu5xeSLGyAcxzDiVirC8cwxES2TkZ1r69tx/1m/a5hf6I3bQRB
uMQia6HWo4lBT60S95N8WAMWt3k5PI3Rb0PCFoe5alwswOAIWSYT2gHqfh3TmQw3Y7tbxdJx/qBi
op4B/izIsDCB6Mt4ucZa+xwazMmhsDWlKBTHJNcquk2IBxd21kLKbs8eBJPORMHrLDDkLEFaE0ZX
D5vdqqu7e9EAw0pwrk5GwYLsq9ElGeEY2pLpkiff2QZcToofbNsePzGhHoSKgNBgn1KW00DnrV0D
19CeXqX23ct1ZRk+so6imuUKDzv3aBGGDD9QoCQKO6aum8PjB9iUrwOfiyGL+GMoG1tD+rX27tOD
imZ/ydiK7uL9MXbkLMXpkdwAbvqiqx2M2eAsbh16T0da/6lzTi1Ukk98nJTDDky9gzwAF6gJ5PUg
I8VzQUgUjrlLz6KAzeJO+GN6MmHn4W8EDgV2ctduDGzE71rdKzD1LZwVRYksUQPSYnRpPhL7Mhnm
Ns/43sMnspEx9VY3fmCYPpt5nzvDwXF2j5RFyrnQ2+Xf/Rbtr79cXl3oC3ddQt/JPa/bnCv9/ti8
mFbEMTlS3Bf2EhDlBefuHRaDklriCOA1Rbx7nqbsx2viMsCBpiONBOlDwUIj7eFrYI7aGDFzV1E4
X9DhxK13hpEsO6YWT2KKS4Ja2sv2J+VPoRNESXE+8nuNOYX61W0cRJq3VBZqFI6IkcjTH4m9Wh79
s/8gUuAcAS4cTxhyRImqmiK6mavBk7w67AdG/jQpTFgHmmF7+mTCOLgGDqoMd833D6/XjrneNNOW
ETNhnFm96agwrHut4AXKCd1++VXTe7nvh21jzbFJL8oDjlheUAmEaDFdd7bzSUs39DhdC9pOvR9Y
p52sMV0bEQFGNSHwgO2jt7DgSdhqRmgFJVnepj1DNKSi0jsThMnujbQow8Mth2GYnHcnZ1DXI4h9
8+11N4XpXw4jecIg5db6WxqiZDaPWZ9SbVaN/qTRYlO6Y3AXAwa7P35KuelczNSKo/Odw8LlGxSr
eeODb8L144JH4Pb8h5o1c38wDCrEZrGHNGg4Nmbqcx0s0grpJ084GsQ5PEZzbd5BZQZuhYfxyqQN
HpoolT0F7mg1xj/2e+kBBe8Jn5a20oG1p7pd4zvenHy1jd6wSyyaaRdu9dp1400kzbWdbd/XnilE
emcWL2+IVUvBEbqWx04OcSVhTa3MnF5eUe48riSVC15PqS2fAUgEgpjG3Vz39J77KrrIrBYNzMNQ
gB9XiRy7Ld8AjHnGQTEOXkOTdz+kUkSVc9y4TE3dgTn3ny38Iqu6b31LJGLOfDPsSmX3Wmm50inB
LkfMLLuD3NWYDavGJYgcc7v4kcm+XgC0BovbuC6k6c9n+dMu2KrgffbZLdoXM1k8jjbKzXLwkz+M
viDsrLPTItDt42M25kuYZESv++o60egdZoNjIyPP4ypLVnMIOHbZ7aJlQJ5p3ci7K9lBkZm6CMb6
NOSkukpisffZuQ0PhVuv7e5T9LXEOfkvbdrKa4lt5tAjJdBWoDKccVZXH5CJmptHzWfzHV3z/5QI
drBAzI/6ILfVhmqr+NRP+IxWzCGhfK5SprJg7gtOzeDkvIUa8/BmtLPLd98bNM4zcws/xj7twgXC
57Ux05Kqg5RDrm+UuySmkvO0LuxCPi2eHPJtVXeMaEfAxvwvVAkUEgFIOjg7htdJbxpvpCiHz7vz
0sbnxvxVlXl8nwSc0ktQmLslvmEfGAjZyu6GX9WL4Fs+zNLh0Fni/ZrH3BRQQKwXnnR9Dxz9EMOb
yVg2hNlY4Pr+kS9ptqfbbuttj7jNdtp1/A6fEyhlLgPSQ8K/9FpA5Zlv2dRIeSyjq74xdYSbTJpt
pmONvpi+av5e4ldBMqDlLnxla+NJUH+G4Da6TwFJY8cQtmFMlpNaiROnLuA4WVo9Da7E2DJB3UWj
vtaguSuzPJMOUc3IseFqfC/mdnn8OjZ9K/nYbnNRQt1kIOE+O1eAVErKaMBqU1qxvAVhyGrKEh0A
14W16/xjBNszKHwDZuvqmJXyB59DoK0lLH1jQN8UZnWe0cRuzJMTzIVrF1xHoMSscnAk5EumTXwP
swDLP0SEy44onXj1UdidEjJ0Fxly3VYc4m13PSMa10nxx5t3RlXHnjv6l3Q+5db59XTdq72YXMhx
Tgnk9+zKoORD+SPS28OvjJ2ZRd3ou7PCiFBwzOPA8qIJdAsYyh5/KrA8303dRATZ76O5HzPKrRQk
dt9DMCl0CiM9ttC9eQVomINF23+PsvRgXXRT0clRTXSEdvxKfU3j7mf3UgO7Rt9p3LpohFmZ6wC2
DzHaYp5cJ7ROJNhHUw7PGs/ZGx8O1PyH1AcxME6ckpWnKAxnzl71VUACdc+8kvMo3QCEYIDThaV1
fdYn2PrCGpLxZuNHNFA9C+foKBhZRSZLel3re6pMq/MSbTJz+95kU/CM4KOjapOlGj0aK3ZNvi8U
ny/W5wcY3b6NFlnoKwPKd8m6/ERCZWI3Y7+TYkDPY9X6gKCmibNyymEEDmF2ldZhgQFsysgtknWz
IRbB4XWq26U6iikeBtRuCG79MqlbohhCwrxkaGXCoVwN57uadt2AY0hRdw+K/4KNXeM1DfKUHftn
4alHTUx90ZQtyDKlrizVxPYQjel/vtsR1RY7zt2ZecTcZ6idLC0tCgmEN7lILsn8GjatO5zCbrmC
gD/9Lbi5K/rdSFRCFQdCeQs9P7xZgGA8KhX/JsFZBdAuJMyQ2+WNctfMeneu+vtvFJBMzXXbef4F
P78cNjzMiyFRUL51kjbvdhMA7Y0xaf+i+ajLvjHSJ9NOupg1ciKewtGBSWbRnptmwVpDalM1Wf0h
otzgEMW/O7m+dEZlWkb8VhOIP5+jEbzJiGdaoBPnwpycftp/ArHc7MjrYjWwfsTFsNcmRHJ5uEnw
teBCXcUjHeXqbxQeeZKtMnM3xzXCKa+dRrnnVdYChgu+bIEGyMtcy+SD6Bh3EYION6+2Jja/j0I+
QSt6dRxuuwJMLJmb/cn1sPjM3+1xEjSBew+xyJzYpb/z0DeJ9KL+2nUxJZs+mhuQ7ajYfby1GTVt
n81XnspQSsiIOSPNgda4P2Z94oFvtqNdJiaFr9JyuUXANVMSHclLmOwNj6YfDqav6D7FzU9sKvaQ
zhS8gU+JQVqA0aCQrtBIPSKAwFZ3PsiVcfjQCIV+10MqeGKft3K6CdMilcP9rTHEQxAUi2yxL450
wCXL2fTlX7QfDDLdvXm+bzhDikL4BHtVWwTvxLtutivt6A7lfzw1X5nGRi0Een2jNjB3K6EjcV+J
AiPbmmexTOzptzYA/NEGlMw/Mo8Nvj/oIEYEqz4rPpJVn11+6eSIh/dD+Dd/uK+Drl1RKiyzMBoC
cMHbirWHr9Inc3Pe/8s+laj9r6A/GBy5Ve9s3bQBq5Jc75pRbo+Nzaa2ufqByKM1Ow05M7bo2djn
awyzJPEBMVi6PcbtFW2l4lkmObMLyejQ6gbXCjMoBvWaHLEelkgq7Zi/z1Au8QeciFNTGEfLDyNi
QjqxctoXPlvcY7dTmnGjCB4cLCbMizBmSd+LGkGJDBllTscOSfFuOjI24eC2FbYayJsx/txk0n6n
keQWXSzua91qsRIP0RtBAb7Hzg11x/k3U/Y3MmY/eye9aznokGZEdbb/uW6Qm59CPo9QQ9XsMKlj
W4am38PG4LdLWeoFBbqCxn6Z+/ypSfCoB4v/kVkSwn0O8HRkI2cUREj+vpLyaUsY+ZnBx8COVzs6
geiPhiRmQmhsKtFaJgfOw98TRFBJjZjXjKWR8W3N2exzCscmHEXqBveWP2N63lEGBm3wYoyeEwxg
vaeeW4Mx1C8BGEgNslMxHWjZtezZf00oNJPOHKQ8jLOLXgyQCk4C93LO/JnOrR/EWFFMg0JDc096
jwUCxj1Ze9kVxZ4DzEAXuY1ZbVpdLBYlQrN14u3o4beH9tvrdUhr7TezmbUKA8FjbpZfFjqJCdep
1xKLYJFMcWEX/98Ry8z+CfZLp1vhe4QAwzLxrFq1WIflzQUkyrsDA6NSsX7aHs96wjvNdZ8Zgp1j
TIzwMlbzpdx2cnqJ6RzrwFYzFE8DawsvHNL98Wf09+VmnkOm9iOgbjX3SJZvJvzwiH3h+gJ4YHn/
xECYscCQCX93eh5j0H0He79CbBLnoiwtSw1JzIl2L9JTXZCG4hMzhVa56+eM+v8ZXJnrisxeQd6d
3yxIfN3rZsMWFhdFnKmolMdLxE9Oo/3AtZI2QTOZog+E+FoAbUAvSbnPgl58GyIztMEjnclQPtUd
tlzVIWIZjUxrjxt+sDqKWDJqxuhH4rie/a46frafibzLkIQpMjHCTIMy9lVLFYA7StZzTAud3dqh
fhf+0m+iEHiH7K1Pgss1RgPifrGDl6+hPAblSuNHc/pWXmleyYlcx+0cYYPVRi2Jz5zK9sfeTTNe
N5H9QmSK9fh2Nx6LUidkuF+OnR4iWKhnK/SymCYHiCQ5HvsoXXW0hMjzmzYlX4LaQ69jshqvc8Zb
FUpBhnIKJxrMoZ3UUYjfdy21kPvngwhlk2h0TJxi/Aj1pNTtwlTjIDoieK//pPOl9ov/5/E8KjUo
x9pHKybUxXKK2x14OvY7wC3+551t51bSSExKNmgj2+/QWJeDOHG+W9vsoivED3UzhrSTN83umYfJ
b6t82WuxR94pFN7biiFC4mJiPdkR5tiG3r7QBwTt4V7UWO6KGp2RDTu1hJ07GdKI1n+eyFFysWUO
Qal7CogLSRTJsi1sFvV8/JZURe0AGR9icNlFE1uTR5r+BWsH8N5NhGnkTW/XOYKMUHkIYZjJGihm
w/WgVT1rJd1OmWqfauyZo9jzcPxAQ2t95z6ITXXaev6PS2yZXEpoVkRgLQDPUiPaGhmlAn4bK5y7
lpLLXbVOMFzq7nukyF6gB1AStyEDf3NVpqoLD7o/wfk4Dpj5WwoAiGEfKtms35LmRuMVEPBL5vtg
SZX42KUyCcE7NkuuPbdGRLt/amQiEQ/4HGsxDssFQNxsPm3fsWo71WdgQDULO2I0/baXXuPEyMoS
fvSuNZFE/M5NAWFY1z+/pRlB3adb7dNUFdF2W6yhANpXyTctqWoqp/ypZvTyQIxnLb1x/hKEO99r
oI+jnjH5rWmCKNuPOBgpJLfq/y89/HZA01yZF+nhOG1Dw+Oh/IJ4IlVVq425/EL4TNEJ5k0abKAB
TurtooV66H6DkV1xGOs+v54t2vLV5ywyTsEWiQaa74E2xAaDyR9vwb9sbPvK69JsS41+wD9plFNZ
B8JoLJl9gdNcz0ADnl+YQxlX63ycM5gN1WVlLgWTYg0i27l6Z5KDLRIrOxnI45fCyPYyjdh64xXh
dqb9aQgM/DOLTlJqSWNkZSdu5bfy9+N78he/ZknpOzVb2hj3vdP2aXFO+fVVjOrh43y0AUyJxU5+
m9SQu3nhXJ5GFO/LvHyoIrjqx5PMTOokIthRv6YDmloQtNtkz1ljuwABOf0lbcmz0Z2cXOyKMqO2
o5Y/zQJDgUa4Z3rCPmaLE8VCLUkF5QHEz+t4E1+5zC8nvtV+hhtXGpSTCgU0qj3RaFxjA5HPq4S5
GbduiX3XgEKjQkLI7Xu0zyHfdOqSvSmWubASaN1eYhZMG65NrTthJ3qw+4q8bzrM8sVy4p1Ivd+5
rpNx6DZvAE9gnfX6FC/n9uh1UxT0ka4uIVTSU4mhpYwmDZ6zs/ZWDvaPBi/SDch7EqmUQI7ICmC4
gR/L41+dSPq/j3kgzCmaaOwBhPfD1UdJlmMtueaEAmDD9meYkt1lmtH7iq27WrUrs0FewdOOXMhy
Wr79htAjF2MC6bIDvrtrtGNotI7gzNHxDrNLg/XJOxM3yGWaKtC8/68B2P+uXShx794LnN5cyT4O
yAklIxV/5F8jU5TDWCxiUawwolWYzD2KmLO5TTT4fxcmkPUX+dscUsU+hFyfOK91L9eejjv1CTUQ
MHeI+VFCpvHbie8wN9ixaY/kmb6JCiW+TjXrRJ4mGLrfM8jEmWI52PueD0o6u750EnzsTNC/xPZW
9cLsPxkez2ea9M6PnYdPe9vgDkEcUrJ9AJoSJaNqME/C/HDXvaRTy9aDTkYc+ODbbfiPSJDWWP5h
9ffOJLrg4XLH6SdJCuxzN0ScPc4EFdSA6L3cO1bgLpvBl/RBZaNsFBpQI2yeF8p7GE7J0hfw0oUR
m48wjjVAGoSyU7ZOfAge/9QQJExhB6U27UDc7O+F1JWhQoqXl9eDSngCFn8w/6TTiMpmp2liuvvd
8m8JI8kVD07t9acRH7Nl5X32wmihfwpfdYskilcJIb/Ff5D+ttr/4CZ1iJK9q2ikZnM4/jlqM7hW
h6e+PDJdQiKRFUUuWcoy+0cgYk5zayaunFfoztdwE/86x088HmqgebcfpjfMagjRRTAezrCR8TeR
8u/VwPTp38fNH4/uobK+lnVYCYGWuyxGqHk1RyfrgpoVxtudsKFnfqQyout8rQzJ9kTJBHjNgjbX
R2btCFkUJzdrfjkU8oIuGQbcfhel+IYAPMwik2Byl77DUb0UUbM709+iPakqw7Eu4sAys8RQItsT
PBObuxr2x5p+PymKU2Fat9mc3Zww0uYE7cAjwL1t/NQ8nC4h3N3480GJolPrDE61V+QcBOwkmZtZ
pQdgklbXEZsb24+ZA64Nx+4v8hlV2bH5u0DC3hMeC63ilI/FI7nzJxeBgA15yrvWOfOjWIxJRjll
mFXNFR1QRi/PhvgcIFmH6RiDeX2DD5oPupsfDcIe+E73RJq0AV0whgrsBGNUoLN9m7fMFSF7taSu
MP+ov7KfSoLgKdgdM6bxHEPV561vHOUD50jPTVHxIY+rxKxwyTXQDzoIDpNyjsGWYctv5ijDVQ05
NARPeZT3MMwiVKc9ho2G5wsLHxOidpZv31qImSiNSldiTKy7oo3W16Zv7yFUdI8z5G57odW6D2D5
w20Zoljlqk6wlHDjPRMtdSi5gOrpJ6J3TXagyDP2IPg5N493+BrgGztlyj20Sec8r7CnroXJ9ZXQ
S/bh/n0Ud929tTGoSREsfvOu2bFt/55dPW9K5a5u8JnPWGEUixq0VsxivmCtU7+TeHkhSqgj+w4d
Oe+wQLIgwjAGufU5LI4fk5XV3faQZE6tA1P1K6/+8vg8s+Pp2rFN94IkeDBxvM6NUBOG3uLpKJCx
23Hrhqg2adVHXD6VuaqovrWxDYnZYIbkSKsj6YiOcLJiOl5aWTwoNj7UKHScWjUPbdn3Qp82cO69
fBkzVFR0dnfAUmgZ1ckgtuNYmNdQe6fiK8IqtxvSrS1xk5ENTdZMnrkvPFtw21me8yVxrOXvY7bx
1iSnvF/qMP16HhVSDu6V4WPV64IA1tmQ5+sOY1XFtUfotPnodH++2ZzQCAfoDDSRiYOaPaGhPi61
Xu+Qvqx+81LSFZN59kfgtCY3CCaE7Jim06AmCgPwqWPgHj6gvRb8fNtpIDanNl+Isv5Y7ni6GCsW
xVEazQCimBHavoOr1J7fJsVejmbfycMo9OwFRE18x6WHWp3vrxqhAp6l/5jD5y/ZJR7BuiXcAp5G
9rOa4VRfzIVK8RCvmun9m+YYE4/dLEZ43f9XzBcBXKsm1waGiV/J0a1gSq+ti31gm1DvjwShIi7W
YKE/hX9W4Ijo3GsjjMA/qQ0clDPG+u63tM0NRNk4tWKhvwqh6o0mYBWy0BAVJLmiZQQQT6qOLt6C
7BRdC+R4/lMcqHHEWDoggtwBrj6Fls6c7NY81thSZmX1AbOfzGgKzfn2dGiKBIHGhtRpQqKgg8ya
mHqEsS/r+d2BsFdf8C1zVvtbeIQZ3xT8K7IVE4+C56j0V4hgTPoq06JeocnnA/VIK9Ur8YwBAqI7
MMLM1okNiAUBuv3arNp6X+mxvHD1Dao2wOP26Dro1EftLRGJNqT25QsUDcj/xq5BkUMd5L1SUkiW
YBanILnmXhN2kv/DkjzDyGXBZXTo5Iet9rvCjAQuMzrfmftVx5o6SpfJec2ap4ARlbO8mN03Zkgl
lEPwpeXxbIi24noMWQbMyry5zmM5WN3VGb27g3Lu1uVp7MUMXjXawO5LqII1ycc1wGFo25FTMFHM
q6sHRbypCw4OQ8qO4IaV39nGVJB5hyP0uBTwJo3UsiLiuMYIheBZmiYzht8PBaIztNzuqep/u6Uu
nN+tfz0FTOHRQwNybbsisk17rH201OQG91Z/UJybaN/PjoI6nFp8SnFGZvxP0Qa/B70zYAwErvYt
xUtJLujXcLxHgyQqge4Ms0/VLcUJZZgEXepUuDdDSa7AsGc2AtOXN+Qto8zBkZODG3qoikkfoaWd
lg5rRmiZhjH6YjgfkQSFsV3EktILZA0TdoMF4Ohc/oOwt4jFCI9eGcflC0dbXJ+v6GnpUgKPnRMP
LtcliXW1N1bCP6oq5BoZmPwGjvKzxi9+dLRFh+zMyVYDkl+Cksh4/xQbrjLd/ORUi3FgnTjKxQLC
UNs7jMU3/tTqjejB4MYQ0DcvgwIfa70XLlFq5vcZIDhS6EcuCCz0C+e38xSlcWyhkyIV7FW6eXeC
AODajGtFr3UuzJscBBbKKD/YjNGps2wXcGbp4W2y3NBqewjNCI1zFOb8Xtf83OPLy4tRAMiaObCF
O4CC44uup7xTksaNuFRcs+7hTXiWJjw7SX+54333R2TeXSHa3yUqbhBC+WEYPtVnChPdtdGitWfL
Bns4Vz2/bM4VVMMVdsEhXfVMlcn7BAxCLig6lnVJkTb0gbiyNEze8bPtrhf3ioE3vxBI8btlfza3
EJqKaFCdG2gwb/irPRZg1wCYHb/Xk2NxcsSNrAEtD/Q/kHPd1aGaj/sYlWu7oD7mN/CCYnjYyDt5
WS/Uy14COBHMKBly+XrMR8AxyXwiovbgXsn6hWhFn7lon3hk6zVEm8UpFawCQFfQd+FaEYOCdKMA
PfYbGdT8egfcG5gdxRPj08GjpqT1wF0YZSELw4sJmZofIZd7o3doxrMuVFhdqzPnXeKibGbtBewT
NNbMrNchh2fFkxeoklMmduaHPHufD9KuuCZavahjW4bGOxO7bmXyiWHqXzPY3sdP+bbVbZ1eX4YX
gLuAuwM1s59+RrR2zwmFaqDhjdWDeTGWN6cPjR962oZsa3PY0ZKznQ1JKh7NxRoWOuQLbsskRob/
g+COAZIroQKnn6rKbyGvbgdgWudGqH6BbezCVntfFsnxwUSm7eVSS+EUtsifySnMrgi/egvZiPwk
Of6EG2Jjs91Q02sqiNgETfs/sR/YQIcwCb2c+/g6JxhyENTq5jk5RsDYcer3ZF+kYnqWd8Vt/KXr
dpOYlLJBK9g2boJxYSzIdMo3YnVWtiPbf68BEeSRWdah+yYSuCivNUG8jgqe6dTuA3j2kkAw2zyY
Eyi5c8JAvQlShfsaGHkLa2fbgQI+BmykntQI5pUT7TlPMiM+XmMdMfx/hKBGC4Jq3FRcrMfzmZ6L
1ehU1hOAKeP49QyBfSSnU3KjfaPgE8EDp+3k4Hn07gBDdDx6JbsrQ7YQHm6FoPeM7fMCnrDWHINL
9MJHloaWUYM5CuQwocBoEfbD7XvsMInQPp0s5ZMXXmj7N90KxFy9W4gk1oSrNPxaqQtMExAeCoga
GpoNorG/rXdigO0cimhErgumwYe67u6wL9CpaJjSJS956/biwEb44OT+iPbyav46HrrgRLhJM2d4
mAhy2bbLP5gymhUcRaLEN1IsB3w/C/XrOrxoArFPcipD4NVX/CI22uw6tDbYTMa/+MJwsifixVgB
/j0yQiJI2oiDNEOxeVm0Pm90MvnUptLzh27Ulii4inKV7Z3Bo/vW/wF0Zbvl6nACJgueJc7dRFbK
IHBBGr1uKLIcPscPLuxDkiyjL3sIaj7eQtM5ra80UGIyIMQ3GSVsaY2bTSzEMcLtfBR7v2UMZGvH
cB827Q4FnXmz5ZsO1dSSGlypEFSEn3luto6bQg6yCWZEsiwAU//HfeGWgg7xENqAfHuk3/81QG9n
vFjxgBITHg2RpZfrWt7A4efAKnWdRx7czada4ihZE0nxTSYewxSNSIwXXkQu/1Yw3tSPEKzGktZ0
GwTrBvCsTHfcDVqU+dDoKlIfvdHU3j9smJ/+YR5LSR1bfW/fDd1P5GTJceXWUApKFMH3Xo8sKQzF
uzgIFVpT2OjHkOKLD8JpZxvyvpbBgFOzvE7rMEJl6GoM1zBW0vfXxPPA9FGl0lvmxev0NhwfrHdu
K6dDJMe67+NI7CqqQhJEW6orr8coQS4yVQERbrZW9Tx02nV7knYRnTHjTBBAZm+ed+BjYziJJo1U
v0oGTNPxaGp1MOXU/hl8/wCOOuF2noG5v9pWrxnGjov/u+k1Vm8VG+JLJk+XAEDojsX86t5oUnnR
X9mXSyL2nAZR/XSbblIaCt/vHbBaRERuVWxBx/HO/VS/uNE0lEACSb2RNS4smBUZTKXvW5oZ89Mu
w/2z652lWt/sHkmYQyah70hy6pzYVIGdhtD2vSRLK8ThpbezQx2GEfItl6Av4gbXEolaU0nULI7a
7N1aWLnsmj6LdfuBm9Wlv3fxXywTyKas7d4s3Zzzk07zzQe4mghwvRjIvKGpPdczCdvLVNBC3mro
xSwTSCE5nMHNpGEqY1bME29UiFPjJjBjnN99KGLhQNnvXkcXZG/jiUbxTyi1CrZfSJ2/BPu4anIY
/fwmGBvWiGaPFyKhnftaNJerfQzhpw2p3nVcQCuvRIdYyPweEyoNII4B9Q9M/GUcgkqnUPYaqZmd
lJ9eK5G4QBXnbAPjmKnhKHyDkmng6OODtdXWgutNUj2/YvH1vtA5AlxP6f7W56ygJPICvJvaYUV6
zjkJ1UhkRnpb+kA0umfVo55jTjd3PVLSrByBw2SouJClGOUp4ROBNJDJyA17sfZM6jXfulOLN3S7
W8eOOKZ1L8I6WqguwIwzNBHN0CFUMyMycl2gWbBd3wU5FhJq66RGgTbQn/fSVKFIE18aZkI7QPwq
PjhJV+tGL4+I11yf+uoauugmgI82553wkYZ11v3/gqO6b8Enkctx0LTy69edXOfhDTIocKzpaslK
eGjwomXLHgotrZ2Fa0Y7EmGtJzyiDwlRIbc+fE9FlrtMrpnlecGCQ3xxuXcSaGRsSr9xF1PB5jjq
S3bcBgW06mdabpOIP5yp9ayTUtjIPab+24UNK8iS6E7Erqc3//ht98NQYL6u21yYGkckFjlsaV+7
FkD6Bz4JpS3qcHb8Sj9m416K+AUl1xx/AqGuP+gCBDh2y58Mypd0ZSXY05CooYilq15VOstCjxuH
2IWGfjQEUwiTFiE0RkLGI66vVhOU5oFRBi/ckPKuUVdF5L7g4NngiEl9JjwUmOf145STLt3AO8EQ
DB1/IQHyoGeEro8Op1qGAzixibwCzRx0oPn9Riu48zEKz0juA4krkTx+Mb72soirCbmJz9L8nbse
3XStMmk/pAX43Z91BBAF8Bfb93bSRmu4Vcf5qCWBW6pPzsXHgA6YwAFarkdKlvbR4X8cv+ISMEiS
K3f4Wm9USKFxzGYbcmYo+YsT//rzEOYbcEKqOnPvs/4xAMisWqB52oTCTbdHKSRo/dpcKwSYbEw8
+YwwRuOTvGu+iiMdtfZswm8nJossvACRW6EEcxLadMEz2vU1WLXzr5OVCMcP+R6DSN5WBvbGU9/c
dtzMHWr5tn3fJmniUDHilm0RO0t5tNu9lxFnsGadI4h6oPDs55RBAucbYIA4q4h2Ya7U9mJKaegr
nzlZSwl7jELW/AysL7pldBRPlH6wzcTFlPtZ5MYYSvmv2UxNVC5teo9MS0V/g5UhybngO2O9zxwL
ezL6EHoh7F9lHKxvHUp4dju6EI+WEfO7g/hdScPMnNItWN3cJrH3VL4jFk4EcvBY/3o+VrRXq9hj
3ze4aTEKMWGBKx/m4TBlFkgSyxmZfT6lpHPRqFw20eFYOQBP5xIsmhjTs7geAXA/2OhkDWfMdfpE
KllF8W9dgHYJb9dV8YC16ADo6vvCeMIt6Qs4ZHdSn5PgOGYZa1m79UfRnlhJwX0eJm/SADatf0Uv
Zvg2iE1UwGj0trSEMGm6R09r2KAAXrVw672ujEqxSpZSTSlSkiWPN0mJ9enz+EjOpL7yHJRkl0ms
PbK748u9vLb3NQtLEkF1InDGyrHzcrYbcAX+cbeAgn179VF4/bb7zDWKLG7StzxgXAP0/i+77aRP
qweaDLCUwJZ9xXfgzbhCLwY8TOMlEA8STKrx+Tuueif+rNGgH8LNfIAr/t9j0gKZG9NGnNLOLGPA
2kRL/yIEDvVWdlggNBwoyeA7RL5CrEQ/z5tcq7Cy/Qn8PxJ95B9UhvDwpaJrwnP34Bl0pPnVAGys
yuk5oMBeffJFFwKOFi0yBXMkaRjMVw7jc2eCsfKF4s5118AhxPI1J8LpjudRUt59cscJh/HkQsv3
Z4o0EiR03Lzx+x/0OIpCAKluu3kOAKAQ3q1+7QsL6efe+sK5caXmci44Oy/RPE1G/Yr/OjwaKvBr
02HoO4PPEoQ3i5J21eXLzxbQVF8D2KDgmkVEIReAALw3OAe2Uff3dKbZyh2ta08+RIuXBzqHDxOc
IIFqbn8wyXuuWk2tXxRRiK9fQ7oc7RdT90chtBCZgpVv3kMoLBXtSkMXm25mkl2pgTCXnGvj+kQE
xRXcAxNzPhzuVDSFQAa13EgtyC72Q2wJa3k5SJvQBeDQLJGlb6G0rimAYzyk8Urti/iolP8WtLKT
EjViOsUVGyEguDBwgZEYOGJWciFZA8j62HZIBMdnaUB5KqRqn/g7uCYy6u/vaCC8KNOaVcCiXhM+
HkQijuQakm8jhofN9iYRwCubfNqKnxdWVWLCgT9g68S6UGTDvGdlk1q3QkMtKDOCjuMTq5MwDPEP
EYPFMGDo+MPTVPAMiOtrnyF5qNOAQgM1BpTnNHN29hIBQLsDhlUypXJeiHwekgkjMHfu8ICsMbSF
Ouy2oX3NjYjzPK1n1U2MpOMQ26a1og7i87LFeApn4nIv0u89OSdEbX84B49PpYfiTQHt1zMtd0B6
GbH5t3TieFXaC0anCRIENw3fXJ5hr0i5HWgfKp0748xws5F6ayWr+uTZrpgcvqB22mJoyqMcebJG
FqFP9lk1GbEENPfRqOuI/KkE4fTD9LTTPfsElx7HccAhQxcBRQ3uM1t+bt6VNFyvRX7jzOSEqULH
qdkrp60IhA001sVsZ04auwbGyPO3X5xMXv06H/bL2nCi2YlP7z7fYPnrz8EnV7VSmAkhl9roKJOB
WDzke8Cse0N7SEdRo1+y/WWVYAyoNMDxCnRPZ9AgTM0+Wb6fcmDVKi/O/XMiIIP7e0No4FRMtFUS
EtpYhdbsYfLxZwVw4jA5YNwJzmPHkBSFefInope4DZrdRO5wXCeWPwKpzw2Z1ZRMg8WaZHayXNLu
Aq14r7/dZdbzK9gXsRwGWL9i8WCt3VjtpMwO9fdYgFqDFE0PHyqOdV0aloGCcQDZNYexsMVCGalv
B7MaQYl2BwBz+I/A7qxs7DM/L2Ml/MNkkaIhPC5BQyEfhqyRrFzcPbr1kysMTSpY57UCLEmwHCjj
/D6hjTYgkHneBVW8F27YRXm8ZgH7PLshZQquYlGwhL8wgJAGZs7XLJ5012y2cCPhtxXG8or1toaR
qpiLaF8F5kFF0CReOptugNBy5LqhawIsxysXEz+9iQQ/zhafeamVZSJHEwuFdMWLokDm7T1ofQsu
ZT8UZ2/Omi5CvLKD3BlpyycOjh6VWnok10CqdEFwRAbXIAiPfahgmST6mkG7xklkcZsNpYtRuP5K
SGsSjS0QCvGWuYEft6Dj9Fjece8VNEKRXzOpJv/hhJnlubNwO5lvuMqjHGjwUxTyABzKSDW/4Is6
mP9nwWXjaVDQS4bP8mGcT8wfbqDljbEtNqlb1f1+UEyQhPMMsnFshUMn5DtZIO89gnH37WpXgLcB
LsfJxM1mp5a6HZdq8hxFVastDKEN0cs6W29o1Z86Ts7JR8ThgjKxrt7ENLSeJD0/3SGa+GTeuJuE
wru9u2jVFMuKVdoykw3LwQBKyEc1J9kBhG+1PNHfNl/59xXUGUPfLq03VtoNGZaUG/Nnzo2v4f4b
4Wo6Tyoy4Luq61QwoXS76AcC45VPCLER6JhqE1lFyQfFuHGxH9mbD0w6d8N0FSylqTKb7DgRWisZ
FiDsTL8V2l3hqr6x2gDbJt4/luWDyu5OlC+YoWWsl8IorM38fM7nRAoAmu9mw5loPzpSTwSozEHt
gS5h50gPZZlEvaIbexUnqKK6WHfr41c3BAORA5elJi4SdJBLq+ei7cAIkdAO/ruL4h3ASUYzBFI4
MQT4ajnqeDvp/JgMWyJa7ub2qFoTebDZGFHkvgVK5mpFTqZbiCOhlVqyFC/pvp6eFfLrXT/Sl2cV
t4hvfmP6GXOLAi8+D7QVumvqDLVifFoD+k5vIdvwsezMSwiyGsQMn/BlmCE40P+ZIw4mhxNFGvkC
9whwIXmTCadu5C8ZzaWJTEvX17+y/mTdZNLfGGXQs9K8Bh0FsihwxjJytjysXxKOtIYIGfa1B1ie
z10B+QuE0rVXUUvlQEygU3z9DIYNrwwqCY02J1EcoXmjtibzI1wLxtavQBaAYc6rHGbRzXahxr8g
rWlQEyBQy96ENLCXHZafMpWq9GEtLkPo04/EaEUW6KKgsxWtPXhCFYVKfokWqPeC/K84hTOmJGiZ
goF15MP7xEe4Ko8HnuMtArNz5cG9wHfuho1S7DLkPNF6Bc27q/+lAQDEWEiTnqzFZ+cnQBlO/Hsf
T2RKAy5tbYCDYX4LJOqQy9nkUEDWMUl7Qrke+eiBgr7LP5K85EoLIpAZn3Mv891vI6v6oztzpC/W
YsO5uBrse4AUsuu7af0pZvxmWGW2LUwqCU4aJi79A+MRWxm5uEzzYG9N5ySEOzjwSWcE5oHJmQHm
eWj+PAHgJ2KrHKE00i4RvEozodvN9uiNT8GFpXv/v/AU29EWJoCsyPoKRt0I1oX2U/6Nx/4hOVdx
m6KvR4U26LIElc7vrv3S5H7L+KmtcYH2MenjoJfrY5PKCRrcSxKKsnxRAB5LGUrcJAnNAIhz4iP3
S21YgzjRJ2qiy+Kilme2PgOZBRsm/1h2Z4+2ZflotepiG93wknC8pyUzRflTzY42n0boqnop7Y9a
5PVRHJK2WzWNmIkq5BWqnk4Cn5lnibjtb79hjnUzRppIgKJOE2ENfwUCnPWF9S50hJ5WiFHaA148
bXi1FXtqsYyk7QitrFY0xvBAIqW3AvmVeT1jSyaTsg9kE4OnWj7sMOdjFXPl612NFxwYGB7iI+Y9
+8Zph/6ePwGHgEUX6ztYjZWVbBRd1X7VATgd5BHhLeY1E7BlF3wjPAtqMMQL2nAGTf9v+tdgl8Cj
sxQj83TR4iIRx0wBct03QiNeIvALIGCd55DwGWrurKBs9181qwNFw80wuZzgy1Fw12FCI4gSO/xw
y4KHdTzK4+61K4LOXfxR9zKC6mTOluf+4iTe/qL/kx07sGvcAjgewaa+6r60sAoPQrbYz7/fDGkn
xmvZVM7a1P4+aX7m4xYkICfVkdmleBeHtWITa6O0UR94FI8+ICc9y5K1VTzKvYkBNg6RqmLXdl5n
VMHDo66CVqM/X/HML71gqBAq1/M9WLpSw+cIZ2auiOIl12Jpb1GKKNRpPU8HiHhxEXnOkB2CKVSO
qW3nW2vkivAV9Ldz79iA7SU/eT6xEowPdSh88Hi4Fp1YALq0S5Udg9It3qaMxClFe8IS0ShtpKcI
RWa7Ptrb/VhLWvtBSC2Knj8BFyMVqIZ8w0Pw9LKqCRYMwhqE5pWrOZYeEhWWAVRTG9V07lMc3DNh
2GS0EplAdIcFy8Tr2XTmYfOByBhbFU2yA+ijBbVTCsVGgpPwfcSJTXdBxjeiicpWJmkYv6ZUGYUS
wm2P3tFnid4cwwekynQZH/ebLO4xQ9lbpkPDrqna0ngN1cqYsnoQdpM1fbALxEs4EkX5RpziBd5B
nrYfgOULePx8W7YrFvVl9FkbhDTMt3/3mDKcfmuX3osACVmuBzl9+/dKH+lgKFquM4hBBdehb4PQ
Z150sVcfoDaXX1f3syCCk8VVkLneWRNrjKqThZT4mAk+YOgkSv8VZdY0zC7PJa5gMs9ap/H2F2kD
ekGy8lTGb9jcrf+iUSR34BwhzTppKAbbDxwNa57ZPHkzWrb9t8LzHrYo3Q2/RwPmh7BNL+08TjT1
J5bXObcwrm3haUOl6tRTQcD0lgorcALFU5b5+s079Y0BM6A/96uITaet6d1pD2A+YfVgMPVANw+R
aMDIZgmXOz2h7cbFtlhsEf+OtW4PwL+IKpVUiacpemxdR77x9dqV3y8C29Z0xVeFVkUsc2z5Vsdf
vvhCpxTlKIsnp54Ctxj3EovpbbIs+4sbLhiTEZQ05qf4BXDWB6kkIqA1rqjftNyc9mIasDVdXDc7
LA8H6rUz/0duv0adClHkZVAYWrcrACTmu9y/WFFzcbMtSxG6PMPN2b4EsAEL89EJidFrgD1T9Ixg
LFMsrMLFtlEf9XROI+KKxME/KSagILqA4DrxoATbbZBj3h/ig1iYul3wC6QHXaA1QveQasOjwB0J
KMkGF73dLdrVfwuwOteTrcWkYi5UpWK+75eL33Bg/1qqJhP8mJDR/294Y3WFI9yBp4r9MkrN1Lhs
evtkqWBUv5IyD/y/c+aEMrWhwFzf9SIoRMgMP2oNDfa0/IYHhJvwzjdNUHBhQRKKPWiAzTkYFeV7
8WlgYhL2FFPp1gzgRicwE7V6LZpoV5vreuE5D+y2L0EOs1mnaMOXnhkfBmQ3LCFRSCpZd6lu88fm
+yTDrc1HM5z7ASjMZwXlXc7vUUE3Op5M+wtPJ3Kv4wYyho5LY8Deoycn9CLfqr1MRo+oKkYt7aIa
gGpYZpoNsfEgDrWfHLuf6/9QKY6/fu8eL0RIYz3qk3GxUhrS1Bc/3M7IRJHKcjQzgPKW+IM4NX2F
Pm3HPNCNabQvwO9j/l7+WQTaD3pszA6PnrFFZ4shoIToEZQAsu3fS8cBACY0IVRUHsnteVa+nOxt
fQhqMhDfkdp15DxJoKiknZYfQoPj2SUb3K7xu0wghxa6uODzYFnWIyb4pkdlQ+YwTs4sUUb26vJy
pCAAmKmmhFiJzGxo1h9pqdd1MXv+puIqOoLeJRaCYeoPPLa2hRE3IQ1GuOGWJX7xAh/XqkaSafPJ
LhEUTTZ4qxBHnnUU0ldeIi10EuI/jJxoG86pm9qHRWk2rXo+l4XmYeEG1HLEwnm0AYEk2nwIW8uk
A9RNf8vjc0f2z5nmxIWqJGJq17GGrS0HjyLPaYuAHF38J/r5/QTgnheJtRNbsWP4dIM5vzMWefSz
lgYkPKg0E0xRttucqQRe3O3hpGNw5r4C8aBBvWfss+F4eXvz0mHwxRgqTYzMx+7674dCUieGawzp
wgbaoVk89ppO8bikeKX92P7fNBQULqjAplg8A7sKMB9fAeBo+iGu8s2TGw0gLp8QeqT8R9zSjooU
FlueuhCsQqnXwsqRn0JGAnJwpjx057WcyFp+8nvtgXLbiK4Ps5z30phF+H/KuJcWS1yC0Tse2VZa
W2jRWfhAoHNVRae3CIeKvGUTcJzlXNfGAPKBO2SdV6N6oY+Yz4zWDIeNPbkmwHNA4lYRPKyHjlBq
0cMVIYCTwjpZhhZLbqXKSNLtxUN2jP68UMXPbnEg/JtL6k8FLcpnbWexKaspQDUHqEx0EE17XdDc
FxGE+BYSlddoCEPMl/0Vcl4xnc2diNKCaKy3LSDtgiLr4UAMNy4vXxqoagxxgYhI9AZGIZsjXFlK
VrVTRBSgMCqm1tx1W0re9XLieI1KHuDgZGseagZZAgEXG6CvnVsziGAU7Fz9OJwlTW4xV9brjarO
twZ3UXcKe/96vYDuWVCHVBL6fJ+QVrR7vYJYwPnRsofa9+/jjM43v7gXjbRa6Q2uMFA/aSHRHxeX
JrGyloQxW9SfnIZMLd53QdXGj9UPH0JOb4gz5tD6RPWSGjwJvH5eW0hk3UDP0F2QMkqTelfWD0sz
uKsRbCma1lUiUYBOCF6ieWeWV5zKl4+rqfLXoVHU0Uam8wFSHVHrN2PpdnvizB9PE9C4UqfyGajw
SbR2gsRjM1AcUfRGpw1ppgwezX8/p7nTjoWFApFX8vMpptkZVPiyMPxwHYfmrWn+LByLu62Nuh8O
GdGfTDwV0izvPUxZ8lEnv15dHkzRGp4ZD+F6FEw9IzKv5nwlOq3Fr0CdXBqZ2nZIIi7/hoD7HTmw
VZYDxxu6ZwQ8rMod6+Llo+2HEgjTZE8OXE6cXZCMYkpEUeq49zQwj6kVJsoew7VOmA/7oQfVb38c
IC0s1iHmeaIp0RWmhqhFkfNlmTsYmTraZCq8Un/1qzi4qQT70T8BzOnntrG11MIqklWmIMocz0+2
1PDj+gCukPvOgrq8pAjlZMQ8grnuFu5hmfiaUcc3pKwg1OxmLODGsLMbDrtsdgxARiQBVQwcyNAY
2X6nvyMY5GtU8L9lY2meE5AHcVabne3EKK18RRPPOMB/7S9C7QmP8n4jDWNfUgd81CoKqCKRSDNk
73dDq1wwaJdRHGT9sgXEB2PRvjlfBIW1A8OSiq2Q/MODlmQkN+edSv60sokOOZDytlGZbIVTv+jN
eNFDDzz8J+lnpSd5gGeURNRFgEizwKm/7uQn3/4Q4SWq10ywn5/Qed1sTsth2fhcKWgVsKMvQjo5
uxDg6HOpfWA80zUCAan3m1PbkULUOWgY52/w88nb75KECEopyH/A7DcveYpZA4TuGEFMJgv+A56T
TMkPoV/FXrHdSXiq2grvnEiuCgH6TLxQeK/HKYo9cyWYU84NMpLph9amYhJMO4QUllKDgF9R83s7
ofUBllBnucKC28ss9MbQliuiEtJ59WlejLejSYG/aTPGTDYhH1hBUrjiagpGMNAxmnF5W2Jzm7aa
414lzKYgJufut/l23IwoOIKADzpqjka4xHVFSVv4DQFvbAUf+6DvbINf1Ih8s6aUeQ+SIfH/9sUO
OTdwF8H6N8mZ4u8gwDdHrEOpqS5LhF6AUlrACYu1e4fi7XUtzOMUSkA7Z4+co4CEKFabBpR4/g1d
7qHGdXbf4veHCf5MneKX3a1U5IGQG0QTo1uPr/HCdkkhauOyTbIjI1rve7Fg10ua/LVnsDMJzdVs
lz6Sf0movsD9tGDKyZWMFUYhDhAs+s7UxtYlwEkBACzXulWLCJOEY4kb8o8b6eBPd9jsCp6xuAt0
J4WB6XhRvYpl+ZxrpMGyOnagQAa+T3+qNXqLnv6YOSKHRKsD4/DRfFC8B2Yo+i791jtbKcZpbsMm
IB1AppFmL6Mzyb+KXmuZhQ+APMkxfmCg+KpAMUdyJCN5KwA+n9fEK9AED2XWtk857wduwJ2/Evyr
Pbpc+qfrP3gTJdQzhqgJwgwSL/WO7ViysC10izqcXMzBrr2/w0tXmX74IEihl3UnncGbph3e/Zam
hK3xBvOx8A/GxOF5xUmOlwHo+PSAHnNXWWEqUVnfRJoPs4kKPOLL2io44M5FBVfgIGanTcInST5k
zxGzW+ieZjDP33BR7AICjVQKfEIjO6e3HVPtQVqv8z424xZlqSL9drYcXT29jyK5W4khfQ4z0kHv
UKLOpuVvOw2C73iUbTYChy2GJqafuCQTKUIYMfzOLK96KEYUThumlwgzHQ6Km/mqtgCX4BjqVhaD
pdSOC/LlLYLA0qTWrBGSxla7Ykhut2Ou0po9eR1Cnv5Q3HtON7auzvK3LBkfycEgcy5W/4ITz+Xw
OazZ7gEo22WhShlLnKmSTgXOMcACERBMj45wTUWILQkED8NRmU5RMvEAmgqBz/1Xwd68I0u0LD2m
sgzX6ziG57Rr0QRynnWrNZCrz7LL+0tyg/6AZZkdunwMxt/Jr7ku6JR0mytuYMv64/1M/pXy8Ghw
GbrtQ9v7XEUZou9RpgqCrTbsX8cqCG3KLSWMBziGDjtRA8sIFG9+MM39xsCk8Di9NL9FlLoKs2eW
NjkcthyCqQoLHKLJuA1vcMpXlWH3OV8mEY2rAR5NJf0bKxe+BAiXb3dDfpWQXljgJTA+l22IkZws
IjCBDz8kfMsJybZi4eT5B76PxbQhqp1WzLwS8aH1IZx5yZlT1PagasjKA3DR5xajqVlIsrrZLZX/
jjm8N/O6ZapaS2KLqKDsnABjj1uVMJj5q7sQ/gcdG82EORfcO1k8bMSFfJEczETutW8Dom5PyeS8
ScKa1uET4dLjlvTj/Ar2T4cCeWvzhFivns0FQ/5bscx3On1bA9Li42EdRjfcr6zM6jTU/W+zQKI7
1oRIpU2ZqxrS5M03TBGO2LOh98rdYShxuYLhnM/m+uayHcTS6zvuXye4TTaAWk5Wxq1woEhd802y
WEluh8XAaxupaRgirw2VIVr8vggOS5C6/d+oQlwmMtmco350SlIW2HFjB4bNX4YIjuV5Ge/QGQej
ye6xcsvrhI33mMbyw8j3HThYNWINxfpt+NQdFAa2MdIER8rvanuJWYlQwkBmn2kIHrWW+pIrHEix
R6nMzFAT469NZXBw0v9t+W43wCVcnOaFyExUwOsTP1TUmBB8iKN//1zyAaFZMiUIuJLv/S+x1zu8
NhA+N1J6+ty3Awc77Om3UgLnhShwkaUywh2V9hwpJa8zw+i2iyt2HkFGuS3wf+/enL9GjzYxOpmv
5B6JJrp/uBz8bwHSlcKMxD4BAXPxxuEnsxz2hQ1NV655zY1O43B9AqW5kiy1PRpSeY18U7zIvHfr
IlH0hQzQOn+MK7cDKEwgKyVWxfKhCZeuD8ilXnJLmfZNJNuRR18kf8d957Qon9oOLoO1w50lXlSw
qFPj2l4BDe/sB0PewwbM65vHr+VRhqw6ad85bhTJlLetKRiaSJmwO1gRHNrHknAs9bFfZLAknF6A
YHjvKXHhANoRa/T/tvGztOwA3ox1GRlMbPaX+k3HKGBYNQFTTWvo9wlt5XGwa3E0JksH5xNN1JuP
2vW7k7QGAKbQNyM2Gq8S9XOKeiEtBFPylgitX9yeVhA8f969BwRTMkcrq9dqidfbMFK2qLVrG0oh
ZiH3cQTlDb0iiwFa5qgm8Tp7kDtGUSU6lRxo1u0BI3whpXID7YQzCwix4MLnpBgH37HdzVBmrP8L
N8wYfzg4d6LYmlqKBonSRenImIA39S4JOgVf2oBt5/M8gVO9pf5sW5s/3nEL6B6ZZ33YBCbQ1D1M
I4tqmqNREbb0fJMGudFF3ctnnmMQ5VvgWqrbQvlfavZYqHAww8tctFJe5FG32xTiYNGx9O7BAFYY
UCUT3PCKIq9E+P7F3c2ZYGFDNsStt0Jd6X+8FF9RnS5iXA8Q4dK1OjOQOfDENshMjECZhGJpoEc3
6PPw2rDZZfW2ZD6Rw1/Iw+QsmNR31sWwGL/gC62iZpM2mClIjV8RClTuOothJegFFArrrD05KW6Q
fNTWaqYXWFtQWTEJ8rolmuqviEQkrvcNoeo6uik4QFdFVdlgYdGPzrt+F+OEjF7fcbiZ4nF0xnti
KFpICw/bWUyBacLlGra/6MGwEB8SYAhUziTrNi/f9GNfqQXgfakGQC/FqhAnLuZ+MhIvieI5ny1K
FPj+zjqwaEUOM177kAiBpxeUqiZcp0p9ELC7uaXivuQ/Ea2v6z90K7quL+a3wS4ywtopTd92D+vW
I9tmAHwbFnTZLGjQA3MaptTMWMUp4r0fefDbWaQ6z7FWoKwsCNW3z80OkBLsRy8yf52nKP8dSR3Q
Ygam8gZ9sWrQgOGJfY/hsynxVnkrBoEFK5qFPGye1XOvqACJaPINw599D+LdOsI9MDKr5nQI667m
khQKpG/YJJk6yyoFBsy3rXaDefj3vDvmlXJn5P5qkVwLLUKymhaLceJh4eoYWQROML3GwT9N9Ak3
gDGIWqoA60N5yBEd86qe8XXSZapEHpb8N9Ep0GL56+KyXbSPqEhQQIQScTHOJKciGAACd4wlb+7C
xzVsdVSqCTb5i3p/QCxEb1soWflfYdrSVk7HGqJYoi4bKcz0JK6xdQIELp0PIxpIYs6oL+Hp4jpW
P6DYw8r4jCyzEkwUZ+7dt+Ep+KV0izrUfHrQIyYa+m7D8ET8LzZVBjlj7Hz+ye1ob57V57NKpL/E
h8un+K3VXPPQLW/eequeDbwpd/bFKcUsUfuc+eGbcBOjrKDvg50kS+P2Aj7fTawZZ4HJZacnhrgG
fqcFc80dwGJZS0b62sWuTf485xh/uoprdVI8wP1c0/UUvDwTQeVAIcBbWKyxPPiZ0tJSr7nfEB7C
GbRkpQcxkQRVlhURg6GX/Ejz0BwqjEmEd2xFlFeWeRMJVsRs9wWQ1v4otxwtF9sxva5nIOb0RTzE
Wta5f9Wb89+pYtXd/SjFjLUagEnlI9zm8obYlk5KNYgNnf9rkBcpbDEGupJWXFoak2iwsM7OO8AX
9RvO0K0mbq0n5PhGDdhYlHEzW2mI1PiPyatKfwKxxE+bHnbfqvB2FINrtYSkWuxKF6r7n2a843s+
XPgBnEGb27qZvbKWHOXAmDYOeCI4q5Rcdl5epaUXzinkAnCIaCGj6xetCPCTywOTIEvCtJSBJTZ6
AeHRRYaTvUrGYYRBVYiD8jzjkUA+K1xFUzhpVxGvNcAFNlqc+AVdoTojOaFecDh2ei1Xig5SL82+
wWBzE2H6QH61roTc43bdybyeJRzXsAanPJnoZrKB8DuJkaGRFKJ8zch96q4UNKkvrJis98WvWX6V
AMoQVTHoyXiI6fNJoV4sU36MTmyZ8h4ETGiHs6sl+ENgIEJRvB5S+7IjA77cUol5OsFIVzr7eEH4
jrvdIGYhbu9fdd0Pf/QagE0nc/mpATLrAtaZGKgNmYCxPMblTrisBYjFMOsJPtVCRWKsQcjLSXRA
OMgCtIN5Z3Wd1vUxmdCZYbHyEmV4h5Kq6BuOSmAhzisrmAw/cmCJXBVy7EinIxiwendtaeq1x8hh
CluyDrrWLV1NzXC+eM2A0bPvbUYMvsPm4tbfaAiCHghUTY6T7rt+pIhqFcUU4oZlLajw2cAmMqUX
ot8WGQo8uCXc1wgFq+pl5NAdLMs6/k51+UHiJZrN/IQo9clyR9zGKusZ2FlYP1v4panQRCX5ICEB
6Qf0fe+W62LBJ/LAXXzsGhgZyc1kynvHb99PWE9HoXchOn8CSXzjeZwebNH3EZbOe1eaWOwbEs9W
GIjxkHOmBHSXxeQmRn62RUZo6IinY1O7YZs1Uw0eskylYE7QxXdcxd0+f4/Xm7081VbkIUCvVOGb
cE0b96YX8+61Cl7+yeLrut4oPwdSadDcsNsOfyoO4TunQ/vywssgYmyczGtkda+JJNNEWKy3az4q
8xR69YbjaPYf+XSdcXyJV1VmyPrN/pb5WQYROPh97xX9nbjXgJg52h8Y85OOBTAd68GEGLXCLImq
xQCdBs1afHZ89j4Pi0iPy8iCo7J6cdChzrkwuTmgg7fePdmSDG5kHnP4dPM95wxaN7m2qfvSs3oa
yiYUrh68MfxTVDI3Fd30Wg/yhvjPOhegwTiHsOgT0ByCuCRkr2AKpwa4HXmziMZK5qXbVh/r0ord
dUaqj08SFV4gnx771tMdc7uX205SXsS7iahGTy3Fld4+bmSVyMZbaVe3eFSXWXf/VTWTVtefecSV
80qfcPA9f+/Q1jI6cg9mZFy8QGvGfHLJNJ9OQBtCTc78x3n2hbzIwy/kcdbgiUNBb4LPmPQh80Z1
jP8/ftwJ3JnbLz/MmqKGHUHg4yhcUEObKqaeaXxnSFvE1C8WasAdvIamZ1Eu4g8ZZJVVxyCh+fJ+
VYik4iBmJIR1WQlkNuYYIBLtLrJZaojGkKUluI4UOMsyDFATWX9++VysW61a4FFX7vwGWVMF3F+s
TNsGnfqncuHgxx32gFZX/oHwXMgNYWfUJIkeA1m9s30cv/bG7sEzfZDmmpKoGUTwVuP9lviCBxVa
9PzBmdpplMNc8I+zzhJ6W5QQ8rzp5+NF3hrJ1yxqzy0jGx6NhBCzM1MfpItBrDEIvCfGuoKdZuw7
vw89X3mAwidKGsaRuSSq62cN+PLEsF+d9fThwgEd09vctT9rvssyWTKz2R+j4Ama7yLNKwYcGMqi
NtwsxaxfJesyXiC75Xg7xg1en72Ct8QkyFQSMvLPhJy5Hnrr9so3aChAEE32lXpDdAY9ZPa34BZD
hNXacjQQ3bG5d8um0JF2ZkePWuXnw/WztoeYtbMaMQ+lytd5LET6HO3gIsqd0eGFDabomGvpoGgC
Sq9yc4SdFSuHqWqGaJTGqp3XqTlD6fuiGNa9XB8Xl+lnB5/xEppfCirbapSIzOjkdIN5Dl6pJOuc
oVn+umf6Uefq7oodWSQ4QPFCftcs4uF1suCCBdTHEh1AfY8z8PD4s7xEfSXuCP8nhrfYCgRg/T0h
w+GVs9YsCH25x4zF3dnThZuSkngCGAe+RWEWFA1QSyNMmkq+z3QtEAny726ctrBzijyGtd5hfPdJ
h4T5ckU/Nr3/fFdC4vrNYdwWBfaHPgv5u0rduU0Vgi4lL87itQZlKX/i87Za5Z9BnRzw08fGCZ/F
2njdvMPbpY8l+eLSVTSb/IbZKcEextZ62IlOUPHMqKWE1eI4h10/oSEBJOA2bIHXevFpiXD7QGoi
7s6qBeDzSQnyjHg6Bjm9WXU1B9V08wVaDFg2+4cuhpb6NkMBAocCYdm4FJ5OYQLv3zpAHeBU7S46
u8EVVgIQ2CwGGJbegVPUnz056GN4LWHQDHGOioTclPWV86POR/Kv0+msMHHWdTjj97fKSVtZDsBp
tCmbVx0//qiDRs/e4fIM/FAvjpm/DJJXMgbJ0rscy/Zo8B/2aDM9lQOyxyearo18BdyyOmBfDdGP
Pmb42Rgd7J+n8xxi3HvaCk2Hc9uyEF1PgbVxSglYStLx983ojjPiqILKn4YU4HIo66HMAVrdjSHG
hLZp+/tsnueMk4J5W+iTh7GI/Gr12FG35Cal7KSu2O01aAfkvbrUvb/4FkMeoNe4PeR5psVJXo+a
E5deG0jZQ6LbnKNWojNMRu33KC+H7kcfi9fdbdz5MmFjjCj/lkkNHwycWvcydaKpZKISAO4tSjfO
HXGhrAYaYpLlQ/zzHAnWMRWAXwiK5LYHT0ukmDgfCXAg/62R2bGjuK/R8GNFc8pNjRohcWGCa9pi
GqIPA/WeEEXx7glbZJrQuMl5hTo4Ohaw/Wsk6/qVuPmT7NT4VCQ3LpLY90ARle5XFQUEKv8pLn7k
bx2j8R9DOfvvA2UuatXgqsUr5ZXrWiHCW3pdTPSpcj1JHRKpOoURS3mLUt+HhYY0q66+n2jmAyjY
3wlsvwAmDgXtznCIM/7RhD0Mh2Y7ZANDWh8B6bhdmpbCEdt1dDHrdJmUS9fVbhjJW6gO8SKFci+e
/PBQXiYE8eBXpngEeAFhLmflEGMcpXnwuZcqENkBuwO5A6H7pBFnBELWRSSUFcM9BYa+icW1wA6l
/WZpbGYPVvMbugiksupx0vnGY0+P5x2yUCMltaW6UstFflWtpZiJ+Du1hBqodHlsLKRYEwrRo9s3
p7CW7T9xPp8e+W5BMErsQjz93/kxbX8dck62ySLUJD4H/zgUdrUx6KcHMFweCc5AuXdaj6FNA+s4
oTurjIQmJCKAS8AxDVrAlp9BUQSlnDI776hLdGWykx2JtCk3qEnJNlebM0P5u0Kc0gElUSWC9lWT
4Haq1651bOZ/KCnnlxPOJVRZRNhH2Ti8i5j4K7zQhz9Qkal9SNDzHi1rR9FqB/h9AaAY8Bxb7yT5
k+EsLSUA2d6KbRpNl3i4/W44+4y/uCdUX/k7qGtlR8kBZh6KD+1Y+jnFBRBvpLZ20PLKloJg/H0n
+xFm2G05RyWxVfGqlYvMRzY5FaFY/KLsU83S93cxKaTzXMWunBIKHeY9ymGB1dkCOTtPrKvf5v95
7RLHaWGJtqmI2JGi5Rsbf20VZGSsspjCX3cBE53OU7Ex9SxT0ZXn38lbXAnsQV8IT8N2uvkm6KOf
TKAJvSZQ/qiT0v1MCWWxdURQL2HIRAAUukIOdIIO+bHcQvl6dqOg4oE3HZGLK18OeI2Z430vqyNE
IGMwwA6UlPJDt8lPMut6iziqsBAtgR/GI2E5DvZKLFvOOyL7BQXpHp3oIw5Tnr3o42YCdC8RxzVo
d0TI2/nPl3ofNcmMikiRlg7JtC/2Em0V6YVgO8GNVrM1+VMjpKvd7egFRQJ1tn7ZssBDZth0aWSt
SekPgLMSJVIsPhqXSmIGzwzZFsD/+z5hQ6fLyW7JdA398r+OPLBFTlTpCoVXVg/jALJItfd16PDh
MNYHrxftZuUSjbmpMvRcNbFsfKBmH2lu/lg822cuY9GQ/X6Ib1HUE4Xbll2N5A+wo5RPDKZS3JNm
BVY0h2Lqx+JcaM06uBY4ZKBjxlbVyWZZudgfP1tcKlbyhIBWLGQHOh/RRgu67bOTHydyyU8Zy5ht
opIG8YnRYuymP27D5Uugj1JX2+DzRhnYO2yie5uWSzMhRXuF56qE7wqyLPRIIhi7EIOORcDRhQai
WIJ5YHvNJ+Ag8/DS33ZXYfTUn47D9t9MDKKdJP0WVbjA6Bk9UK9fJEtQH6I3mfw+/nUZ3dWbNeSD
8TEdfezs6rWkj6vjfo6/Xa2gJODMonduCQqf22rxCVpkY0UmcyK5/XLrCgXVWlyQImpl9N2f4tEn
jdN8RjyfeJpZJRDloIRSqOjhjnqimObUGTly8nFgaprrqpFfL2RTO6QOH96N4Vhw5i4D3v0KzFtc
1NNe93f3Wmck9rPOx+OhfnyYZXxcPemYfH/hKjWtiBSPojUDx5nWGPYepsvOkv71/uj78DMI7rCY
hwSYSuPDLebESi+00zT8qP0Zeu/Z0gGMLcwnlQtZ6qWaYie8x7qsOeII3ejCA8zgNRiLPRvLEepO
IR/jr+PwmjUj2NSoQ0S4gYZpH/uM1L+pCmLq0kVJ1DupiS0MZA28yZT2rg+6JN+0cXc7bhgtpdPk
Zm8CbLzyppvNLbdOXAIevelBS9/rN78T8IRwxH+t6FysrzENEUNWjT7PuF691f9hSNTIEyix6ccs
/t1nhVbAXE3OlPgdMV7R0FmwcbRAUQXwbPTM96r3ij8BSmw8nVjcHu96j1N68nc6EjMpK/khxj0i
F1SFkUT9gvpylf1DVIHDwwbtWbINk9YRQhE8Ldgd7vc4/GwOozoz4rxcb9msREQEeWahGzIC3MDo
i1aQsN34MB9Vz+LQjHmLlpaDexAZQBESdAyGXXOWjph69KbSX8QzQI5wyxeOLNhZiiSiqYBqnqAP
M5mF534unIU0XeIrk8/8IfqoOdz4MWDmljyycPsO4V+RYgI5jTLwgMiZL8E1yMzI+RD2HgRG8RvY
IS3YhEX5ZI7e7ifRr55qHZTFcNm9rhz/pdtudG4bTmIH0ZK3XmLGU1Qm7DNR6D/KYSYvtKXKpYAt
mOtbJaCCg5LzxZUJMLZ9zQV9zBHPIi0GfgUmKq8ROlLn33jh1IMLra1+NT/BeOG0ZijQ225cfFsR
nMTE1mJE55dASEiq81MbmUjcS9KzE+gSQZN57TTk2bIXpkwHxunuqulDy7mVOvE9oQMJ7fiek6fN
0pdOVWINKW0KKHXob2qO97iazpSMBPqaBpTSRGkV1UohVcEvTKiAEvgnPw9TfFaZXrSfgRsl6TJC
X69fk/Kw7VJZ1FB40hnwFh02+yfWn6kfgx9gxvrAk7hnoNhmLTeGEwysB4yffTZvwG8vfBzx8aRx
hx35CLSkG00JYLsp7j8sNH3s5ZKCCFiPMl6oz7aBciPK2WkPHVciOl1L23gCjiT+CuWmBYli48XU
WKaACHxK2juECJUT7b/g1xFc0aVDj9WlDqbwsdIfv5fRyniRDrY4ashxzlXXJ0FU/NVIguuV56ER
7amhg75QW+qKdGdIhSZBI0PXCc+X5Ijm1nOdn0s0pYLaXq5X2RuYtIYe/IYBn1hy/0MLtiqxpZPq
ccDw5bOkr5BIIOk5zRHw3HrKNQSOXnNIRWQicUgn6CTSwmO2q9YIn/8hRMNUvjNJIcRNf3G0r3Qc
mm6P7oHwOs7GiD/GjrQy2RsxBPN2/quXM6k9YJA/3/f9MaMbAirQKAhQferYRi3Z/urDrA56YSh1
NBKytGIGvR5HIwOdKyLQMoSJty1JMlpFpuflWFWkB0n0bf6Fw2CT5wFW3jiS5N843mQB5qjmPWzW
bKD9TbbnghaUhcypiw8GPuIwQaRsXVSmuCwF68GKuFSdCDh38CWavg/p3Dvld26qeTo1D0U3oZou
wJB7cb+eazdsueuppLw30W+RUGcrvlBmNRHIs8XjLZIPgM46o9zg17Lwa4U/OiCzd39z3I1nnDfV
duGdSxY0WepMbYbszW6dg52ttZk9iwLHPxO+YDmO2SWLTVSlHrh6TxpShrWwSiFsk22jHhicyKQC
QiIpDZDDudmyIgRoaOiVedfXPoi4auZtS+oNgBKnCjK+zcJl6JPeuf/1RzhpmYIyxvSwQvQxwfxC
uznnmtovchLIaNPvg2XYWo/xvxdRttoHWHVYwW0F/qxLaepD8WryN5kLVXjtj7CHckS/rY2hZmRe
+cAaZDBpgNNutC74nTjJUt2d24UY/onf9IFLhFk6Do+x1KmA20Nt0dfREzYpxvDydVjKeueMBST5
9wBpOYzyCherE5ZWjYvF5jLxeyOZaKNskEWO4VM37UQ2Wi7JtAms20BChuJYW9wC3R4KfvPEahUl
XoNvG5JG8Cl4fSl/cSVGg3v0QuMAqaJplnU+1UoAQ3UT6uWK7CNW1kByGTN2kWcwh/D59fVVNqgU
064AX1jm/7SNfrdHbaUB+cjxWNe3ud9Nuh17zXMBRaPyZNvKllyzV9ea4wd/ll25QkCV47ilxB3t
MNizOoiupMZ5McDl8ZjFe0nxBRuIIhVpYmhe9s2PalAMqnK+41TjpvD5WWkxeTWj/5xvg/S+f+kF
uZupZ3Li0N/o/8qS9no1tY9rcm+HPDtkCb3yvHLVD9xGsznJ3BySIor7dntnx7Bdzej8uxrP7ozc
t3lJWQPsuZHjJDglx62TLXwxQObMY4Aeb7y5Af3+s/bHPzAqugQtgtkb9KBXT1Rk03SKRqItMzsW
m/lEnBuC2bs/Ozt3UKJuxCf5szYKuvo8XzRzNHEVFiBWUZTB+/YuM6YdcyPAUBunUxrJjq/+j52J
PU/yO5Socx+a33Foydut9HVxC7emM3NETU63zZ0GO1WhtP0yI4m7TH7U4GWFivB1Db/ANiiGhThA
XHWQsjMqeTfVazVAu9wVZj6kJSe2Wg7tcGo5r1ixUF9N7fIv9GchooT5kIh7JLEDgLvacaUVyR2H
uKMUAAF+Vec2ZgxEQVVTJDnwqq2GkSBovTRpbqR3gBzXh0V3cUxIlUCMSK9qUHyIH1oM3uYIp2Sc
chydQJpUi8rpl5hIadlkCSwnCWKWd6m3mo0P9wHr5tYJvSnGQWjHpnfe67TZSxHxJ7q5atYZSu/7
dsTngGY6q+9YB4sTduz9gLql8ltoAXMD/IIrulKxTJDFAeMR6Ix0xYcxt76Dtz1P+VtreXz+uQ3x
8+HKyA0pyw0NHnLKe793/oh0ieAhdgXPB1CL0hS9iFAMCIP2IdHCxWZtzHW6ZSWxuOSaTV/Qr030
oVymrHHNohg2BpZtrWqClH+xDQ3QzjATpgEaPNgolQgccscHWk7H8AvKTfTL0lJiM0c3KwNx34KR
nW8JslK6euEHGp5TvOE21lVhaCcmj9BptVeZ42Qeaf2fvCqIIWOcjmONse2JTelAHpGFgagR7Qcw
Zenh6XCFc4cikEjX1H1smKsKx/o5425vEygnDXi/sWccablT11aluNm91B447FtFj0cDvM08dMJj
QZZ+ph66XodqqdADdW80yelDqCYk4u46wp5liT6pgusAyhzcyzjaH8ud7vcm6yePSCMBrCkV+BPk
kraDIQYq2sG7OCq/aLmkSj40UZ2W9Y9DmHhKjj8p/o5VsfCggrnNWFI/KVEYKjh1lqFtExISDadi
NYjLp8aaiKz1BTkdF7jaBWL5CJ1Thj8w2VIp9VbcmMHpEuRBgiCtLutgwrHFbKrQtUxeAiZAa+Cr
DaXtvZtTKF2vodCdc7jz7S46qDBHpiua0WAhuOudERoUSMSBnKGI/2+OBan3HRcdjzZq+wcnAEmu
RMxQ5n1KQNtezjBwCFjeVcEFt5fbFWI6+vbCd4zFJ2CIiJ5Ynk6AebStujPb/CQe2U9Ql3JTc0eF
d8WYrTzdnkZ92itnlQ1I/+38PhMQztDn8ia29fUsu6eJytsM/EHK1gyujcKsCUfdEo47I0VzW0Hd
qgxGv8y7NlqfMMel3b+8Lyer2h4SzAOATWKAjeuu8MoVew5ARIbwl1jQt+pYcZHvkvDfsuIc64dI
IvWsR6ZPla042ZiE4OYSTvwU61/wlqg8GU6MhNDoGXsrDYefIzLgCyqJ+RxbEuoP4m/FVEjAQzPF
INFwo0XUKy4pytxd7SkA78HlnmyaYqn6rl/ZWtkzVcbnD8pho+bZq1x6d0motgyspOsRNo2rTJ3h
NnwwjKnQp8uFiGDAcSHSQfJkD4NHwTZdnvWvGxy+Ymhfq54eegTh+UTA6ZL/w4R9g8GvCBz8lE+b
Yn+enzI5xOnncrjblzfEpi7hWB3SQFTtELlDO/5/SxMqJgy/zOlRsQCre1/zuWzPQMz5H+4j0IZh
hPK8FLw8vlx2hboYut8GnYCGR/YMxpPH2WPexcOf++iA1MT3XDebF+zw8d/8AQznPdOQdrAdZM+Q
jg9WkluLLcipB6P0fseOmivQcm0Af686JXc62byCg3XTLaW6b3tKgDMCpvn2PXYLJhB0gQHuxwDz
I50cigraivAtiBNnGO9sim6mPmc/HB4ZC2gCZQj48tHSJccwmdMY1+rm+xZpghNwpYT11MAR9cKY
J5Ru3f3c0vy+UKIYJUws99ZpN21cWI4eR9sY788p7aY8RZHcYJLsEwAmHgU+70sh0BC0fUgmvm60
eDQlYDAdCmeiUgHrUGMEGQbnnHnA8iOZ/XvJFmeWVUFW92eDQ9DnLY/D4uvvxN6yv6DLypxR86a2
uBHDANMyTRwX4xY+CBO4GwnLckm4EmqIhyNdqQi6Er3Q9Ov2+sUKF2If9Cqro7sq3Yx/Qao3PoQG
NlK9LXITGTympaigqHNW5N7O4B1m5GTY1UY7u27nTZS2aS0NNZWAGF4m9KhQskAq5z5XWPFQUEwf
hXRmNjhilGsyAT04LHABaGSC0kczPEsYoIS/iEwa1aAXJtIVN/+UqbbQda38GqLcSnc3UCZaIX0B
/aPnTsZj72HiSz3UMrVWJhnSkVGGo2ZHzcl5wat0t4vt9/k9wtNFg/LE8VXC/4tT6/7mOfBWC/K9
/Y8quhK/hUmQPHIsWRCUlcLTbrhq4c0IXAdnMPoPnQGJ//gyEITabbZcO+ZH2jOpUHrCdEz1YCP7
8fAkOI2F9E4+kCGBDBL/lMGZEvdN08dgfr2TxEpHlQQW0EK5k1e/KjtQjpek8Z2/loSjBdgfTI4P
wKAN5Oael68mcB6MrZxfqq6pk2dmnSNEPaXowu2CsYAgpQCHdkEU0n54L3aYixrgnn729d49rqF3
eb7jKy8w8AFpacT6Jwm4VUv0+uhBEIAQrY7//QTxLwt2dVEhv/cQkI7WADL/B42P15LXxyrifXhx
QHBmlpfpZSjtwG5se1mKW195zlKXfnoDfDo+OGm2f1SCklzLh/YO+rrM3/UA85ARSTROn1aCmkCR
+emUg/lRlFapxCPmq7H35rkikjcCI1PsGkwweaykHhIpow7Qshy21nmy7NZbxD6dDHtvq9vwKUF0
D4i6HtHYSyH2GM4yq0bawQLxjMX/zx4/sd9FPLBxXjdEvH7VuOGBK3z99CFoE2iCMaVtPQzyPiu/
+HKqb4PTJho625mBXloXJRaF57jmyvlzztdz+DYWsMnd0XZXa+qt9rSUNIxn3Ppwacshypd3CvRh
9g22lnHjcFTm5i7+KAGkBAwCoUDaZ0zpyTjrcFfY3dXuThbKEWJ2fA5o5ibCkXSSa/BP0VAMzKAN
/9r8kf8r/ctO8RRMj29vjyY5RFC+IMBERJ7GEzvJawtoQiVT+tGVeh1zk1Zxe8l/7sbSga+QESG/
iq3ezXCXERHW63L3n+bOX80AiWgyzQU5A35zPyYY1ocXJbA5/W1X+x6YbiQFB5BRzJ7D3DkL8Xa8
DF2TVZuNc0M2j790KN+/AIDpZRRL6f73YKV5NHzuzovNIySqFzJgRVJGEIOhwj+5usPuEx7jWxpi
JlZadilL0WTg5qfp2rpdo0XztYl0gELWDoR6ZJdM92uBPMrK5PB/1zpX4JRupEsT+YjMZYg/7meH
H/ifgb4vhXzI5pvBg/7E7wg21zFrpStMTuq4W7SLUlf3nneRu/6SUhz1sG7AAa/xI5HBtPlU1Qu7
TzO+WmHOm6xyDPHvE42DBzmCKaULGbhBrtnkXwlpQLEgLxBydo7alChOprGEbD/Fgduc2xFR9gSr
bRME2UH8TvO2vkKn3L+OqGm7HApaVhs+l4gIpYRByjjATqvpK6J/+I+5SDZmu+wpNHAAs12veVpV
1mgH/QMvgeGEqC+oapgs5naTgzNDsj2qvPsOvCUhbCBMWmvbuPxYeInql7AMr9Cifz9NABAHimMg
R8jnE84B0lqPHTjJ5tAnweKgMx7mDoNaoMhzV3D4rczOusAEBBQUogbL70VljGEEmON6yc2NdD41
LdsGkzq7VJi6IW0V4T0HzUt72cHShZkwntOm2s59ugO8Q5z0QqSg10O+8/F+5BDIf8rQlwWesItz
uHcskhWX7pfqlgd8ZGDgteesgGEA+FGTd4GZM6Vx+PYXvDqY41Tq59xCTi7TjQKNHOT+i5gkNhZ4
DJq2pc1hZbX4+mOxPzQMr+zpPV8GmGx5OAYDjIA6ZCZysBhk6H/VPNSt/bihdjsQTb/wVeTesfjd
YLDhQ5NdHGB7gN3Hvw0ji/9GyzxpBO4wHGmR9g+css6yErAhMBDs/HkXlEZQU56EvUra9TMTyASQ
PzBvqO+YXwRYPKNqcL8wXa+wJpHaHNvEQ8Z5O1ed/1A7AUmt0yT5teDZSnQ+1+fUr0VNiXtVCdU6
aU8zm9kokK/G0jFvo4i8BgG7ONnphoaCkpv9m70MoSIpKnswLpRzj+jHYS003FykZtN7nYg6guDQ
vTjLANVXvYpZgNxCTx1RpS+tpaIfOcY+T6kymyQw83R6coccWyeNvPXHuxTmVnDbLaGXHUKLY3/r
/n0JIa/uIizOkW/N3Fe1OUBszYXYoecxtKrBFhpsw3SHyi47jOqkPAxkhhgS1t9XW84ki0fa+nLP
xaEyjMZ39XUceSvespQEL9Qq753CPwNDnTy1x12pg5iEK/PQI5/QdvpSQ48biqyRiREpPHE/LqXP
SM5Ld8hMo1TRhWmvMyAL7iAlCTMGH7RmJamcJrbCMaMDNLdJWswXDuCYh5S/iIHPK2n0890O4f/0
sD/+1ClkPAdlW/aLR1RWuCKd6IyDa8Zlp16am90FiYG8w8GuqEdkjWR88j5jdbMmnXeAM1/w2Y5V
PhBGw/N2oyjEK1ceZe0laNSnVfC3kTDsd+yrAAvGwxs1O2CiTRfq6gA6CkweH7gl3koRlA8T4MG6
svQmCP1CO2fbGTiHZKHy5FQ2OPjkgxGL3CC0tjEO691toYURdwu3PjBWr3be7GlOPQHO55cFpn2w
fsgTNFVqenLQPqHzbkKszndAkST1Rj+XNSJSbkCRdMDh9rt6xW64QgupB/tqE2kJy+LLnAGx+43c
gMGwAoZLkdHJ2spPGuu4F1LTRqTKsPlVK5kQE0s0+fqrXpH26k21jfLSO3VfXVgwc78yQmmD2JbX
RYa7wK8sboeknGrmJL2v35pvAhB/tIhhz0DpZXmEyIZnHvM+QQ8iW2U5PLWmuH65ilQjbTbjtxhw
jQxBOphGKuxAU2bbohA0PdIXLPeltAvzsfpvGgYXS96+FHQf7C7RneJPQvQGjqUIBXgahtoVXUop
mtesSniJHr1qXuMi+72OdK7teR4dHxYIe62/i71nTk85t9jc+ab5qhM/BQbPgyqpeT72oQaUUWLW
CGYSqOMqvlD4EFhRR29lQ6A0xLZZyqcNcqsSupsfXKyBYKo0EkUkFStc5wQIdFSAON5zIQvO6Vq8
V7bvjWqutPBvCXOzZ3hscbG7QcwMhYRQ1tXP0xmO/lHSIqssE6l48ySmsQKWmnUZOAdZJnBMhTtp
/eEW46nG1lYAiMbM6/12Z6SjJyVFTwUi+IafZ8HTmnEJk5GIMccUoGYZRkorUD5V4foiacG2pEYb
jFcLCPGwgnj6P71bgpgT3gROM5ovTJ3FXxOixVjLlpVQhxZ9YQMy435dPdHN3Lvmu7/RWc+qrJyY
EItgcZQNeCNzZA0etrEhXUTmxCJFZlKw03SQIsuJ/Q/gUlGi1QeYoHCPg4omcefDiWaq+R7zf8gd
xo1UmbPAh4X0gFKhPORCkpV73XyMdPpOCwjqg696GMk7h210opWZD/xydxPcfrnHsPPElEXzpdyS
lq7QoPKFXUOOL0uYQVcL1t55RrfX5q6FP8DCL6IQmpYaEZ5lM2UQlU8pslqpdrQYSKWauq098XRx
J9xrYw1D8C9/zKYxRY1p4aoQ2JWwiVFLR6XaOwS+y9jKqk5iMHrxJVACZhxphQmgQOHzwT3fD6vp
lxCXOwI7JtvVEXBON0hkWbMe7sFDmjOQZ/11TODBj1nnzhn5eemEGc8CyJ9oJIJxxzwAw5GfSvxs
SWDD0fOg6hwYUPWq3LdfgdT2U5JtgRj1FJLwbsCzM8gI7RJrY+MdJHRiIq2AGE1LYTlilFvG2wKe
hLj1Ncel+4ZFK8g4d+TvXvIWluxHgiCCqZZ6w+nr/ZK9HaiaL37At7l9g+9u2WqiIw5TBhuG15lR
CZjJcZiZd/+8fFV5li7N0uP1yQDsE3lWj5JRviZGy6EThZEMyL1EXOPmxCBmO31WC8L4JgCJK/9F
HWIa6CuBcLuWOExKx3DtFM8cnkMms3HDtq5Bu0ld5uOojQ+1unIyNeobv1LEz0BEauIrsC0loaMZ
HOR1gVhQTBbQhESEeP9y0QvWLdni3/+XdVncRtL8A1U7lSsC3CyC8YgAccVsUE/GCYDdG866JX/O
4N/ZSODqa92VS9MJiQxjOHpBMlFyqOJnGXMF0rec+kbEacUCpZ7UO6f+RL5fJ+nTRXDws8v7u0Gn
uibxICE4wHeNyeqOY6/6fJVqr3y/dEr/yHBV8s1iIsufCMuqIYpMElGguVB4FIg7VqoJcs2V+eid
guoY3FUYXWI+xE6JoHQRPCpV4/wH/8Mb94Zo7nBlV4oixo2K7Kk84E82gTEuvxxdoOied81JCG0t
vP7lmCcOF4TXcWcrpgI9FC5PI4YZ6AgJ969dQwCPxb0DiTcLQzGYjrRVTNjltzUL1OPjDiKWMOUq
6aq2uV9I8TahTlWx5S3m0iH9UOPK8MmbKyYt4yqV/Y90gYldX5ootmq7CeoNFE2o8+/6ukJJADkP
/U4iBXce99QrfpKwTPJCKCfbuWTkqfWbWGhCgzfHTEI40ZJFsdLpOQ97QZqsE9XN38Wi9RhUGLVv
E4iOmdC+v1rdgwcBI3xtYhm5r8tAEb65Q9bk6dKCrYDv9cdzTVk0G7xCC9vZV3DQrIjx0jVqorbh
trTohvlTT3Z0ISDxBcq3W31ZgcW0tzOjWIXjuoCSrk+vioKpBs9GNlmQVyr/sKvrcqurAm4Z+kLs
hCGS4qkOI6crVG2c2BjbxOV+ZEP7TVdTpPY0DX99UMX4slBBHq48+9AvStr4uOoMWcEom1hzxjbU
K9u1Q5Nin/z7YgLUhTB3w4MG9tBxhoKuZEW5cm27f7YE0uJtlcW3GXLnvvTTK4kJGoPOY4bP4xaU
SkpBotvaP3pKyyD4MBN2vVHQ91jCgDlMLk9WQWOqp9AXgFOUYi8phWTEKw/xfUeZf8AkNfqqamFG
8PF8y1KS1bJPAfvXlltWRis49Jt1KNpAezho6nm73eAP9+dEqgX5nBCyf0cbTtPYX5lPUallRmnl
zbc1tx3ZQzNVFwi2KIKF0b3om7vD7fFZ8ix+GpEDapD0P7m0HWM6uqtBUiLav/0e/4AAnh/XcWmg
8d3Y1EYctjl/zsTgrckLILS9YBXserDhCY+WI6RxNa7QmnCwdV7KDHwrDmyvHy3xtDQ87Py7TZwP
7R4lfk+NK2LDtbP4erHlTaBGW7xCTuoBeWyIUnNkkezXgXSm3a1+y2/LyJfyfAAhIIjaxBzN1V9h
TMVQAM4AkOK+t0zzO/uuHpxWtYJTVPlKqm/FD7GxmI9BfvDP/+7oLbUX9pm/VOA/I/3pGkzRCVd4
sckRHLLmPFAsTLimRWTBPcaIJfRHteLFSl4wZLRJnb8RkwRhlPT/pyyw/3bnb+O96S0K7MeyNkPK
jKB56/E+K0z9WQY3vgjoFB+vJ4dXcgtx0qohVpYQ2tMQilZ4BLrWbgoTrZZ9Eeq8tUPpRwmc1Wo8
pySpQPyjC43LsvC9up8Qctl8i2ojm4w2fGvOIqdm4IKyymTpZlSyPI/ZwEQyhBroV443DEodYRVv
ASybTGsvsS/WbK37hc8gquuRSxSbF1SPyUaqs5Taf9rGOLVGQ5lS5OZCQ8jwCMb9xyjl30h4lgB3
4vW+iD5rV/3g51UgUN9CreuHjTNkfLRnd6Hw9HLJayU2bDq1YRuVU9CzsOtwRUBqCE+fvDVuik98
lO9g3E07iesj+znRAEqdI3sSFKP4+tW1zujjhimPhG9ZUgMaeNFJnV+0aeHTSmbQn3Mi1Fcx77p9
vd9hq0TKK4GQS7ZIs827ZXjjQxNiS1m20OwIaQ8duZBa8YdMOwq4PxCDApjSzTFpQJiHmrPYtAdf
0jbxAR0R7slv4eCam5kfQnNyjDGiGhsdms44h78apKgJ6jFYPR8gfO1FnvpMMmKLzToH7bFFIo0c
HgNsNg+YFXBeDv0eg866MvWNrk7zV2JfQ87d6chmUdLPz1QSUODJI1k6NQrqJaXTQ/XyByqoLH50
3B9q40QgcbkdoQaug+jqctHiKs2hjJPrgWBu2N4C8/XveaFnWuhY99O5Hkljkxtqia+92UL2+3cJ
1RJW06SMoInqDcn6+pnTSimqXu/AQxDNsTfAs+AeRd6RS2+Phyw6y/PfCKfMOdLbirLPTCTnLehl
JDGkj+FlywF6OQb4nVIYKJCM5BEJHVaJPrnJs4NAlCbCUVW3XJ7zDj6LIPKxcnM2fRVW1HNbkmqA
P86t/pDmuBH6tPrZKO2ixA/sQaaKNUXrK+VcqvXbCUmVFRMwIbPowm2Rds7CTqnQAM9+qda7QuZC
wySyNn45+ExjXk3fhy8L+oB1rHXtCT837uRqspnrSD0kCqMrCcnhAqDfgxGQU56TD/EZX30Jnbfn
nOABuuPCh+G9V+IvCy9jLsnGY+xI26uxj7TWSMNQ2Aq/m07jpxDWNqEnUf7ZsJaBe2hRkmegAg2z
nQ6GcBNKb7InSNTtwkCU603ecCoRkfvAxV6bScWf8dgmCu277uUY8KsQvYaTb6wFJVprBbKr7RF7
d6+IoWV+aAQ5rCmjzrEF0SFHEE4tdrFG9NouwLBVdIY2h5giSTzh4AoPPXCllUGj2Y03ti+yegyJ
m9P2J74foGPe79CIFqEHwgmz/RSjTG70EcePz60AL9LdzphuKLMILofbFJTP9x4ULsKjgHKONtTR
fGiGjV98DuwWGHx8U1lpKyQqMjQKFgXDjeSDd+sQuud3O3ZnDU4f28+uRpXISH6B7om/uUY8LoKM
gJ/m12TrI0M0MXvC8gncFkurghkzlfmNhc69IzCGsl00crUBHAWy9zQjxxubqDzzPd7QgBwHsRhj
sEAmvs9MqdG+gyMDV1CT+QjKuyPWlJcu5s8uhzino7cDfN1V/YtMjWGmjL5ULuviIg3vMCgUUcWJ
VcnwKezVKR5ACoaTJlTXknE3AMVX1N9Cz6D09YCyKYpnlGujvWMsyehJhupvkUQmBX3z8oJqKwDP
xJn5RRfPzi2Uic6BkcGhd9slLzV7rcypwdozZJtIdgRkY9Oai1+VyZFyarctVrbCFGmLYcvW8tIG
fODL5oo/WUt7oZlJIkAaggKRNWgmsQOEQyXRtAGzta4wHdItp/NAO9aU7jGknilMjGnW9isz0VTb
ITW3SlWK+hEuHIQZ3ewwQs2T77ent/eghqtVisiGX2qLWnFw10CSCcH4UqtUIX7FOCOar3a1m/8a
UwWK2ED+TtI73DBtTm3tvFtJyHprKlD0UxqXyA77BHBP+QJ5wAXqldKw+Tw/RUjvPqTVy0bQKBoY
rDUN9cbhsBqEPz9tpxxRA/OOUnPvdD7k9uAQ/zvtXd6yToM59TCsLunlH2Z/Gj4qJWJghU6BFi/u
326Nc73vL2AE2SBRLAyS49EhT9odvnM/8JPp6HNIDOZKVZSt2IpCac4iB/I1So0ou0hxiPuF2Hbh
iYOlUjW6h7gtQ/1pghJFRP7fBwQdewfTMmXboHowJjFFaIhbV7AfqmXt52h1VNgESqmrwnu5uYXN
TYLKMvwh5qJFfixN2GyktT+5tBfQChGreQ0ffUdh7QAGJQFojQ1QyG5avdx2XOx59hR2WRFqY4Li
em/rUHUYR5XmLLNN1O6H0mwBAe3Bm8rAVlR+RhBD2XjuUXfZVoQvsyfuJGQZeAJHzqYHBHG3jGaN
2bYh3wreeECiu47n7VYDuZBASF6W3SivN5rta7vSsn/oaaWGyr/L4+zEpZC/2uIdtHJ0lpwi4QCy
LDVGZh1RM47WMfbTeU2EY5z3KKAmJnOC3SCy/QRGog2kw7fC7k+WlNbVpuoWa3J4DU+ltYmS07Gz
JdTuB4/DxakhniENcH/ggGt9M9yG3eOGIJEcB5Rlw7iHpornSWrZmogUeZpXyWrso7kCGhYDgh3S
LJJ7BUukr+xMTGnOUtgO4El8/1/LoTqbq5WsthvIDzyHmXPuVIGxsP3NhTcY/1roktuPqz+3EUKm
GnA6cbI0aTMgKM1UKnB/Ma4ScSFnIxohRCVG0i3M+nllpzS6D5aAO7x1kgvSriv645Mwf1KWj3m0
tqinsC4VZJ7BGwOiuOrMLPJQPXVx5jQ6IVEKruN1OZVhEZOiwxF588fTVS+hivhzBZ2fiUc6wITD
VScU8u8oEbAAvbc/Vipce+OLxGvdx0HxVPAnvNR2UxHM1hHl6tXG2Vl/BH85/UfYwbFOiJX74eRg
8lBkVv3kCE62WJ3u7iPUMvTrnUDvNLK/WPMON3HYtSfydQE/m1vlVvVrJmyqI6ZFHa5rw8xuvys7
Dty6CnE2CEPquGKnuu4kjvgmJ3lt5pnNBn99EJwkX9w2kOcmAl+z7OKDPlh//i8sf0ER1btw24cu
78nOc8atQPdWE33piTag9n8LI13q0qHaaUg9/hG2e05fKLlrtcGHixZ2KidUq0F3iH2vEA48F/M1
9rTy9PhtHz4LiMe1V2bsciSQjHi8+iTmHR14xUk18RdHxlo2V40VrWeD0B/wIrdhrMbBIOMXB1BH
HeFtKEEB3uULyPYPiN7728VH4Hgw/zfS55w/HzbJ1nspTuEiqtSUtdJ4KFVuYR63T1857pSjgF50
ojzZ+eZIp2Iyky2+d8AH74Pjm0FPaqXxa7FmZt9qDOwsuM2Bmp4KITOfNDWiH8/EyZhJubawkNHf
vGvZs0TL3AQPbgBS2Bs3oUGGpx91Y2tvdwBk+JkdzsOS5UGisKnBPuDtHiSZI2v1tDVkYJ421vbd
9RZoES7X+T+Jyuxdk/wJUFsQJU+0RSh0/8Vx+bvSwnIBs2HL5PqGdjJ2cZJhmxyDjeHSNqj+m0ri
qqAeufRxM7ozHdHFcERY7e5yFXjKHtBCZoAz0wP9rzaJiTHKYtiWMljcf2JvJggB+5fxopa4stBy
S5jR48NjW31zt4cvR2MZ7IDORhjO/uCObnsEr9dW9HwMtkwyRCZFdDV1ZVedfe/UGn+lDMdQwy7I
DKLeoXJrhv0DZj0P1oQM/QdLTlJ33gunhtcdIc/8jVR080ksrF5K885Xr9j1wnTG7TP8zsTI95l1
CDlCWUIzrG4kx1PNNyLx7laZHoqwdkt0GUVNXJaUBsBNgP8yJn9p9kaaH44v9+2Sn2TL2IVKWB7/
zs8cGkSSfna56ssLt/FOzQLQAyoESd/VqcFj8QjrS+pyC1RRCGgWsZV85gAQHbBy4Ob5BM5JXIZp
5iCFXSyBkbNCATCzY5xYWgiuLLOoRegoDPFAYOlaHuaHyVhp8niWAl4al1WFUE+k4iKjiuBzjgUr
vocV8fr4OO1LjXhqu1ImE/2cse0iO6UHyKguOkqgxcRIKi7/IkNxFVgUWVSbCQxTSBsb2t367PMK
iNUv+tIJvGFDOslerysyTOaOdgPIDw5qzDtiA6elC+nSmfZ+1MhRTDrBkt0PZltUcVB9fV1GRplf
zb9fLabue4hNtkaAAVB+5Y/qMbf7SF3dK/ROOj6BFxTjKhavXYizV4cJVl3GEpSS2BhQ+j6jVq/W
PG7yXoWaUo68gV8DsrNICzs1oStoLYS8C2PZL9Y7gANXtJd3vNBoTV+2BwpjKmgY+gFoI6eFxpnM
MBh9Lvn5SJQoAg5fYlOkHcIJqvDde/FfyNDKriwjua4eQuFGC2kupLzZX/Da89bCF7WGQ9xk2o6T
icby+3vGcz4O9pXXbXTPqNAIvTBBDd+GZmBBuGuQIJ2Xz76TWvDBVl+fuDXjUrlb4yZqDMvdnxpz
lngmxAh8LmkEUGX9fLCcjJYxMKnBniucoSQc9E2dnp4MXHzvth4GnZgUoUchcK6/vtPOC635MVSj
QpAWKSdjeJGUmJ2JlxlzztpExhsxel6/agj7gMBGlG1vwCw7j2VNXyPgrzY2kh5k1lOX6+0yzkvq
bPnrok7T6Gr30g7GIaDdS8ypNw4n5ZSy8ScRM1NTQccLGdN/6xiPsXPnem0D4msntQMlYLi+eOq8
O1P0OP/3tKtNMmCLepY1MG25YHgDoKGcRJNlUNa6Gm+PxyX4MNS2jDyHG90m1wdMPgbE3Yv3xji4
Z5qRWiTGP1dvOnaco38vZ3gVwTpmGPsGQG95uJ6qBV74gd5uG3Ax03nOHBAPfZOFPyOPH+y0V/nV
as+VXkCFdOza7AoM4axBk1uXpcJSAmjRC2es9HmjVnD27nY4WQsovst1wZC+K4r2vwzSVwRcmQP4
JBqI/XBCrteZdjIe2V7mTahSqP2CCBLid3yTwgAnEGtgYV7wb6YAGN8wOTWIVLW1J7ktYqMM1K5A
2shU17t65KAMqKvYga7T8C3YKtNj+6SHd+cDQU77s7Ws3r+ec0miwzdAL/DDLzufyeIZ5Two0wOI
sc4btnEA0kd2lWjOEQM6bN/z+O4KeggI426JFapt2FstrLDLLLfRAjCM/Ts207weNqYtDGMdbfGY
7vdrU0dqX41g6uJnuMCYDTUInpLCVj+dsE8WcYACJlmtAlljIvqNSPdY53r65Li5PBB8tRZuIC4i
7R2aQS1cc9eULK+d1ENh76zAuNCtwCU+tS8cyEL0ywk0pFs/+pBSIePgnu89Gs1OnG0V5GDGr5zX
qiMAz6CKx3rwjwm8z7t8Fl4LmixSvTNQbW2fJ2IP471VrSlgWZuHnW1NsZa25usXGf4o6Vi5liT6
Spn3cAXjtma4WULvJ2VhIeucEmxE8N/TjVMYSROjo3UpwJdopnzbBycmoyTeyjSfNQhDmOD/Du76
FH4HPa7bF/kVljlfr3B4wAXh83mtcGnZPWuOYi9m+kF3UGM8bCcsj8nkMghoj1EZOdnJnpxo9qPW
QMKTjfvhVSrSdux4i+FJyS5eWFTzd/gOZFixF8W1t7DrNK9t0c/nKDhD06k8cbzUuattRNKk0ryW
XJXBcBoOihRmbI+fEqCUp8EXgO7d3gKXgFnJOgPrwMf4NEZ8Fk0hDfmwgV6OzkjhC1yFlEn2zmgg
z5nSj7v8tTWG6JQESloFmC10rUBSCGl/JDrCyIPcCyzzzKWtGeWk+09cSxGFETbpVq32VRA+BykS
n0AewY3fJ7slyxf/zHd/rlodUFMkbppZxUckAfNZQonuYNrmziGQgbDou6YKUF/hTyujv8v3xHbP
h/hSAHxAdBQZ5Fp6Qarr0IznAwFnHUcwQMKK6cUyeM+OLjnkh8fp9opHZ7vYHfK7J9PfxAmFveY1
ZTukbenKL7Dg1XKQn60bup0HTMrStZ3M0ZCGEFwzh763cHXl8Q2xhWo80Vhb+IT1rfEBRfTprE/x
BlLJmzVapjRJKxbQLAyTkzG1Yo7nfqXgso2dTZpjo6vvW1zgntWElndQq47EZXJHeCPlnhKaG/zb
klzfeEct0hMsqfK+r7D/5moIk6YJnNwKlUQmWRvksGba/1dnAzgYypCG8EWhz3uE2+t1pyZ0OMbX
yTr2lVP3rUvXkPcydtCua5Dsusy59qPg2cmv3H3IDdYgf2+Ime9UtAxqmTqijUwEf7ZzYnhcJ/7D
zUfTlA1zdIf/WUf5wGm88BqLSJ8Wl2eUoo7EvsEuNRWdH/RpPec6SCXRxP2uhTK2uqOdK1oVn3Xp
pQdvCw5009Es5V0hET1yoN4GRkTYZjJg+rG6YY91lheKwmZqbaiv+GNFZOAXEdeRLOiDvLbKJ0L+
GOotVJ9e+DQ5IcgGV8LEldDYPQZghb4J7E0N2B7fx7pMy8U+KSvU269DYXjKnGYWTf9ClRJ/ICBC
gHHP6JVZQbP6b0rwCFJh8fCrqe/oYNhJ26CNtl1MVw+sSUNbMiEcLLOfi3Xf4bHhPMdWregsS2g+
BYJwAo6D11d05nVFohG0tDf3frfxCy+etV3Gz3mjDP6fee3uUYLW0AvBZeGxhfv19yaUQHeHxQ69
j3e0btU3+hGsJNipw2Mt+FGe38lfaZ6fiAw+jNj+GkRW4ecDK8/9BxPLyTRxKnTM41ml3vKsmASf
/PwDQhSKJf79Xk4h6PsH9RqOAupubAVPKBKdFt3Bp3jRRfOLgxzWTYILEbMpdzKCCXynrHlpdJjp
DZ8EC4JfI8V7xoA/wvoOUcjLKsmNpE8CWw2v75q1kzPb9KjPA13IUHXuqbRyNP9aqLXlVqi/qJu2
aYAarqFA3LbiyZhzBy1wXxTBzd82Jl4V2QVOBJwQ/hPvOkgZNd2nbcWp734MGgK+qs6SRbjQUv0v
giru9blBH7L+LhtYYRMnqxaNTaIHnfX+Yo99G98PEFQ6n7j175wHDkrJu0s7OSGdW+25VhGC12MA
WXo0/GnBwLYdFDZroGpAecxHee6XqQOY3JEG1VyfdcXpolrp1PUg5kb583OHLJXzPtsqOF1WwgGu
bHW1ld7Xi+wj3xs4taEE/p/2p4gOu4XAJ9oicGGS3vnJyRFt2SnbBX+aZvLnO1HnPyIRhJvOBxmm
TmSm0mktIYaXYq3qKAJY85N/H2ZC2l9FI5Ziz1pXXDMmQ3xWU4jMjdobVUvBUCOpd+aADtgm7IVL
EuGiF0bsXdUyCY09cVY+spzJkeFbX0YhzuwlJV8wU5cptib33hLfv64h07ekJwRFlmHzVXur6+ww
xOUxxGsKK8+xJEm8fU85uV01NS0H0Mp2kGNhH8lwqcIj2/PnKv8ZuOiZqtkaIesPMQZiFXBH1FiG
UlObr2KIjADv+nenjDPkNakEPUr9K+N9lUH7oUU8Iw0de1F5QKMQookhtYYGNnUlpTpdQZf4l9Lp
NsNnVQ8rtkqme+8+UjiPKXNUyp8xIL6QExhLZQ9BwnM0dfVMRc9Pu7VJYmDm6f6Mbn+EwxPweLB6
HrIsYajLUhSeNQTaBbKWSiyvHn9znFqUmoatUCbj1+lHz9EygJAShR/l88NM9PmlsMMS8byLxfP5
jP7Cuu8E4nHChj2LW51RjVXSaCmigQuaVXvtJ93KYqIHkKNL4eXk1L4s6+x9FqxQdwvzRygXsXyS
PpZgAnkLIvcLcrP83TtQiEpD/nbBUr6LCeJKjVY1SeNWfss05VJ+eLmaMLbwVO0aS8SitAAd738V
rKs+6/BxOQe+fLzqSMEUZhzbONdftShJalnRjj5iRxKaCRMCK3i2PabJ4FbLM6iPmNy1FyoUMN2D
fEvvy/QjHkpIy4glESSAheVl1zTWzmabOnt5sRW3jp54gowYXBujeyoVXAzcYw2ZySxDG1BvRL/x
J9yFmOTLcSh7tXKRXknaG499EkthdLXVW3qkb5wyOyp2MRROcWnK7xegG7vhwQJbhTsrFVvXpz59
/CGC3nfvDMOcwwTB49xll0lc9524i9Jynk62kNi9h4u+l20HW567d4BliGPiL7xpe/lYrMDiPd+N
V4cIwffu0Dowfvai02U0s4puedx3Clz+Uj72WBYDl5+VkU75uHSEdUDV4rIW0PQasPkxQ7gVURbM
tA6WVF/t+drV217kvSl/YLMch/WDLQScp0bfOuMNjH8YwBjFAWAuMPi5IBHM13xq0T/oMpb45R7N
3OO4GVFD5nkPbSzs9n6G2kNSo/tb5Xqzg0q/RtS/jIMRZgFBzRMA5rHhIgbCtpk4NG9B45u1I1he
k82IN0XpHtgk2eWoZRgYSmXETX/aeNnOJInn7v9YrAGOc9MZLNHyjWbf7snodHBlG951IouL4IN3
PNM8yTxN62RdM3RVr04Vg/xeIwhGJM50XQ7uxeymyxjU+Ypp5DieYMAPzd0SHm4lKe62iFDsTyCC
wMEvqs1UFLlwyiX+uCvap0e/1c0ynmFwqmMI3AOicAPkPStUa4JcR/NfeUhAtc1KdfV40wT8dVni
Xs9Hem8erHe/02zVD60zzwfucLE/wmm+9SyfiIG/VcjuXGQTCOSaJ9mogaMa/rLYyt/WJXHf97Jh
+ElDhd6uQCYY13A756TnCxt1FG+KSlN0HJNqV0peUB+rpxituzwzPuY/CvMfkizA3t4WA2pBLY2c
dzzvfpTnWSsirKq8JN7AYwgno8dDllor8pDgnHoh5oe6XMQp/kyBAUE7JVuE4T38tUe70HzP/T1L
q3P0UZvXzjc/NIcfFBvhQuDJ6Qm8u+y6ctIC9m3+LzNDUJoIVJaHmtAoKkeJtuP0KZ4cQphTxhJB
cLzjQhPa19hp2KZDFgH7b8DJxKStqPO4d216sZ+w0IFPszcN1JUsGZlU9CPno732Dt0aoE3Ho597
v+aiJtBbMCi6OXzR9AkgXYfol1se8PfPksp1cxSO94sfmAHErrSdvFCshA3KqmE2foZb78V+mPIg
/+QZju8D3FWoah5m71unlqgyJ+lcYertCPzBkvySfGZETiCNb8Ti/b520cufz3HqxhKld5/kNci6
S1MuM8K1D01W2rcGexXGYURQEyj8vE1/leOAk64xwp3goVWVGd7H6KdkJHkdYDMljliV9KwcAlRg
VPaxptekhbkMkljqL0XqFD2WbbuEciHKkIGU8B4ow8Xykwq+bMsEDVe1DC/xHBE5Ltg21kBGu4qt
tQkEzKQNiHsob1AvXscKqNLT24DPsTbeA1V3NXSLynk282ZeUSY9Be26r49sug83Eifa6v9ZwC3A
4+A9+vzVCkhMqu1Vxo+D66bKxzNOIB/eO379Ii5J1roaMk1IsJnhNgKd7ug+WfGkejAZklLf1d03
Q4w9QDKK1/W/Yv6ewc304AGopOXU0vgWNxPIfM6Qpyn+CCJ78UIHzXwjfZUXP2B3ujxdmSX5Amsb
yVua9kM/HLn6/CUrV5M8jUmjx2s6UcjlBo/0R428osOIiyvCuTuS/pL9zoeEHJkpY7GTFvc5ia/t
iZKb+0uJWNS6+8i0bOXjtBN2Uom8upWhRlYbL6TT3up4eUZhpHKStQK+iLTHgQscLTUJUnBsSd8w
q0bPmolxV0V3aM1PMIETqaC3amhsUn8YZ1lFposrznXZphW+cd+7QCZw8OXB7UIPOh7sD2JCkdd2
P9mhFd9LRySg8XcQ2EQuhVOZ5jTee8bG2zt7kLyFx94vE8FPHdSRuS1LrepAgPwzAqiPFl0TTUGi
x5Ya3meAPEkI0dRLL+U+CSNxgD2hMsOt5OQMWDf7nN3l5NP8K/E6iVaYwW3aq/5KjtCGctjKkjLN
NeC2kDs9Lca74YVCzvZ1sMSEToEjqXIDLzdEFPt8Swe7KYb1O0IIQI0Zne88jg4sp2q3SQOQHtkc
8bOUtemP0REgiLfcgFXeQ1jpUTu991cFgCMHQxTS2csAtB3qbwOe8VM1DJkiY+wekLFOIQ1PmvFu
OY1Q1CsyysitV09VJ1OXbGBc0DCswVwFyQjHne5MxzAJuFbZqLWwmCuuYfbvhCKJSLZlcH6P/VMd
lzvRW9ooSez5Zf8Ftb7nHosBPvoMwN5gTO7WquEEaaCCyBIgLIcxKSncwyn38krjCp8ocEFZtsz3
iZ1Y6aLlJrKtscalqD6n6mr0F1mEuOcKCan3Cnl5Xg9dvV4R4/NexzAz76Phi/qnqfpCyc6yG1GX
C8tIvKZ0scNnP1l39We6eQMxSddGS4txyu4uziht7dfWI8a3YxNf+5wYaBKrPE7i8QbMV62IIXyi
bQre2eHp95A/rMSWEyb2yeFIknvTzRAsL6/xQq7G7lyUuU7WR+a9L8aC2xXVd1HK3zaFeVZXj6Af
alNZZVVlORspZOlyNXVtGFL/YAZj19Izm6Ij9BcVZLiDyIO+OfuvvF00Zn7eTxd97ByWmymcnN8p
6K0UfutNtwGy6mKeqgIr542K9D312FNp9dXfnZnrBRoqHB1Re/7/yvOFGsaKTtUn6w0fG7wRtecQ
HWG6dgwuyVNinzufxR9nr4HFOtU7bczltKSUnq72RQJEsYsOBUvfYrS7eJkTlC2dzHLTs5V8nm0J
MUdLSJOlIYZmtHhTVuuk+BY71Dbi4ABWlfarVfEBk6yS4KBRVV4PNdMta8cjf62hGFQDFYWBB5KO
5/fGy67p8f5O19I/n/j5/wNlHwtTiBYlGu4CJBEENfnBqh+q1LJ49MNaSkwUf8i6Yp45+W1VxhY1
L0szKvuAmRcCpbwj+GecomyjnS2SlQb7gpseT72s7n+8B7nHGUWH1NyFixYULkbHnf1o3+q1X+QM
ppPyYgLGSG6if9cLoHcc/2xMeRsLxhcWGm/iLsCi7fnm212Gh8Evn0QyCuN4XiSziGZBmHoic13l
AuhPaED36zaGJijVovn5UlFmu8m5HkcOaw86XA4WE/fEAIu9VqLQG8RKUv6OBCKTAfHMuIgDQFAH
G+mM30zNk3qU8cyo+qKJndi8HhX9B2d1FssAsaapFoKy9QuRrN3b0lQkZHEV8k7HlI4/jj96zZor
cts8NMGKtjt7H8lAuPnnra/AHaWOhidZcR/zeCD4Z4gdaqoesFqIIVwZBlw6ExOaH58loaDlhlFh
Pp2sJYIsy9Nu235QZtxC8l/1PciyctYDezWPqRkvl4TzmB6Qkp5ysBTilDHwQv+tHS96pPDuU2T1
AfIXpEOO789kKyg4ottAOgD1w7rDanW9BoYQLTX4y/1ZWWRPKNRfqQ47kHxrK3qTvRZP0iZpup69
VuMe3XXy36MeLTbThdvL16Qa0JIMF1PXaXyReBq3y7AJhvc7/tsnb55dOFN3FP14Re/iHhTwI6dd
jDTEjxBBjAC3txZ0ANq4emLoC6qNCaaLhC1KDVf3aEU296qK3OCwY+OcvVKrBrPu/+wiBnQLMcIv
luDZczPJrF2m+lG0uauOvzkXbERi23bRksJ46tabsqjOTGsa7XOr/8jox3Yo5vL/hjH0FOkjMRan
J/p1YtOmtrkk8jip6m28e/enFNlstWAbe5G34E1y+AzyBC4Nth+PTT0zboo98oUF/odw4PMfKPB9
B1QeKu3LLOY2nIjVO4oRu6Xt5sv3DwkXFzm2qEuT7DdzAgSVtE8mgk8QqW1g5ihVeCGI5Iht5TKX
H14xYrEY+6oA6/dV0I2NId6YOzZc2e199JjimI3I4Ell67At6knaNPFCwbOt3jYFJCT91eA6QINb
xSfxR5LVngDXZvSHp5L0l7Ht6IQVfwGriFHmO5sPh/QEh79hNwJo2bXIQEu/7YDT2BSQ6oYO0A28
7rsyv8JzR4NlomrF73KAsmgFX6oW0K42q48Mrd6zWV8+ExhmJUbP+3dtNCviO7FechWjpP745NAy
27EiyRRffMke1uQToDKZQ6Kjc+oTht8dYxDoA1/kHq46fhGdx9y7S4lPsWd6TR49uaBFx0PMb8gd
6rQJCqhTlYEuQ9w0PJqia9Q00kEh9OtFb12zqQEzHI31/2pE3BLaoL/glYbMhGcv+B91hiIsGHJf
iTxtTWwU2+snspMtpwGpYT6tViln/krsXH8q3Wyfj5iQNnU5ILki6rP477ZAzsoQj87cLGR+XaPo
rqltkv/visS1oMg3Qa6q/CZV3T2RaMJqTp47p0rvwxm2Kq+CzJg0lVaZoKibGGRP0p3CziYgSdk+
IXbg0dlQPiN+DnTWPfdKxg8hz3t10UrGdfx3Y3S4t6NCfbVXNzH9OokVbThhmnTsfijDHZRmIc3q
7pRPTuScq6AUmeFXVsO6+zV7bAa6uWytIVaeHIm3y/N/nBhQOxWN7xZyPQyGT0EEjTF2VXZk8WA5
Dplfl4XKqA1elpHBdfI7XWiUuORahpbGfPovD1GkJsGroWgZLpmp1/itMsgPnY6hs8KL/RONPQk+
u1iwR3HKRO3B62eTLaSsKqLal0mHSPpXEpTTLP7WYzjTDr2BxX6Fku/q8c06e3x3rmJj+IFo0Q/x
PSjSlMVN088wHM9eR48oVxxlh6SmiYfnJLu/AuVc9FE/vxfhYCVjQXjXujAczIwMjT4uHUDzIg1u
t6ad+/s1W1dWiXGeCpXrjquKYcyVFGXjzjsUMAZIz42yEHLFtFA3qtijCeNR6u0TZNDHhHbwBsOG
cSwfrfJW/XpPKFLz8O5FR0tNVezZ6YtmU+hq4jELQ038wD0k9I249jLAHUlaxP1GdE7ROw9gR0jT
a6FkQT6AxDYmWe046U5JCiWMN/0SjkcoKscGeVOGZzm4pI/JgcJvFE5PLK59sKqJ+GkjpbHSFPJH
KkDqqpDCKKlykGqsqCrjF5Ij7hHenktGH4E5xCtDrQVcRBpjBxwBfuYG/cCPJcZELu1m4B3DLPAs
xsl9POyvGDUqUTXMVBEmBLqnM6bN5/nV24WnzRarx0JoFkDcpEBB4MX/KjhhG5dAJt+Grn00tzTD
4ovEpwha7SXgd0pwJjygCdVpITT5t1Kc5zBefVZ9lwh0Oi8fdFkJw7+NlsP/Ik7bwmueZZqO34jV
QhSRwW/yNFV7fwb9lkF+AXRFh0cmZXyfeDS8FIqaRQrD/RwidPHmTzP0/171fHXhVzjWGmSgtgAi
MRcii7DvHYYAXNuZQp9EA0L+kY6gzFt03gVwbrTcNoOPaLucyhCsvYRrTlgdhmf7I6rBGts8G0dz
o8a9+WRCoFgqG6kWRqm6A1TV/yVKZUqO9jCCqUYuAvs1Y3aFhUxo4Q3nHDJqzIqPsSqXp2j4XsLh
cn48t+FQPwU3Witcj7eCACLQAgT1U6e0vlhbrBvVw0WZN6MI4Sbc2uBKnHkIMO0Fk2bzcLm/t1sz
uJNHegPBOorirp8CBsy7AYLGH/6v7PgszcMPIh+SyXjLpRMZdkl6PxUKR/gkiOQpxq9HnFudF3Xj
0QUG9DI5L2UN7gWH0aIUpEGaOJSIuSSaGCtsNAq638OVT/fzwcje58XY7gMbv3f18oKke7iNJC5P
QfFchSyiIE8Nxn/g+DH5zQneXhIQV2MZ1Xud8ILGnfc6UCgQ8R3e7xZgV5YjZisEvnRAM4teqzdX
cXTT/0Tgc4w2s9AadueiM1E2CRuxAv8jFZRTQvgXb/wNRa4ySHq+L98jeI0ci7oxBkbnGxGv6P9L
JIAQiTAOvj/L6+S1V3hhqxLbziPQEfNnHg+BjV9f8c56Na97b2tgCAQmrQtzf48GwYoCx4ARVobx
XhIVC927PKbS0RCcYXnwzLn5MIuBk+HGQEWVzd6m/2Hkba739kkeYoXCT4+ym+4USTjj/+iQ0YRR
TAmvS/W+t9UIyJNU1wBqLQxaRVQZRKS1ZTBjn7wTihxZvBIJn+DRk0vxIZ0wqfueWRXV/GYc2h8k
up0OOZft7iAGnNkOqKxJ/9AQBmhAMgaObpNbkMuyoojrh12bdWwHH05rf3lGAcXK+dgkEiSjnALH
WPJWsxxaRcmLszc5kWJKwXKmj2l4isxEhFgcKEO/qj18wcCoK0C2PUAqy/R78VtGxtLrHh/ZF6hu
tX8E9YemmQLRa/KdAAIhB2EqRbly8ghdVNMgK5yu681wBpBcSDgUhJ76a/aHzYHnIBc45/OqLusP
9Gj7AxjXf69/d4DHPzYC+oMlDqRd8u+C9Q2dyalxo3OJGMk/CNetMfNFdHyWEriAZIudkHPvSfIr
5OOGQIuVhXS0nYGiFLEY+1oA3jSpne+ftGshpGflkcvEl1P1hdVosAwQNvcg6C8+LLJ08VuCFzYJ
9a01bkGqt8ERe63MGU18Ku5UGNCYX/d+2WV/Ta9Ldn8GwUsTZqY+XrqAbAYTbvuNda3MPdEtrT5Q
FUftZ0TQjQcWStmLZ3STQTIMTud0R8ZqKZ6JkeVw0ToSzXK6irdavwC3ooa0dNZMFm32rN9qBy35
es2t80Wec+VXiqpmzhYZ+QKtcA7xBTxnkeCX1s3qExwAi3SXDMLpb/Rt1R3bebkHG3uegfVb7xay
gbvKHQrpPJByT8MO5zkQUiRaBQrOMAJ3tpm+wPUfxACaeUJIGpTIIpsnz14VfX+IjaMiLnYub2Po
khb4vYo8KVoiFLS9YdFqu2+JbIpDErnFwqyHGJnlpVa9YHhpUaQ9fF6ywnznpfM6Cx6SYyMqabza
C6fd7o7y4JFDg2dftF2N6PCDU0254Zu+rare2AVk9QRFetXEgoSJ5Ow7/W1jbz6G96VFuNog62cK
6ZBTG7Aza3xyuuGIIOwsTu8IfoP4aL4ia3rFImHe+XsJMYqUWuU9jQSutCdODNqzMJ1dg+Q7xquR
UnVQTbs6roRGuDdq0sw8jSV3/jXLVuSovf2WtCxrfxgOB4DYWmPNv/PnDtZ806C9PtDHu14Y1mxK
VICdtIS1rcB3OIQDUc6gw4U9OvgY1iLla9cAguJaC1871YLxmV5OOEpLKy3aCkjfRwML2F9n5fsd
s6JsPlnWa8komllZs50TN7btRV9SLgn5m/bnxCRpjdwIzR9tQhWbrcd2zhaHEtsbHc1ZesOp1jyN
STqVSHHvFoFH93saLn+mUyf3dz97GN3+ErJgjuYx1yDPPMUl2X7H/4fWRFrctW4zuzbzbpMLY3+c
gnIxiN2Pv7ie62TZNZu8ibMgQQPkL5bxPSKMgdTSyCGeM0fCErQcGa4FYveCmktvfPwX+oWWTZtl
yhrSjIbk/rpYmy+XDWSEhRNgt+a961mjhvDME5eBtMX/D5g/DJjQlpksfcYGmlmmDSZIt1VFIMUF
XeiIdhro3PeSr3sZ5Gx1oZ30kQhWMZZN2VCfxSjxTA+yS3xn9WnWCNbxkEGHhdqLT0XbqCz0Oba9
SkeRmCjPW7SsO7ag5nGHQL8k7DLIHSouJvuwXWdGH6aoqs16QNWDvJOhbFi9qzV+OM/LsFcuubnc
YIZe
`protect end_protected
