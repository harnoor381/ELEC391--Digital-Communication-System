��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����,�1	�)��&��(��H����dP7ɨ���:��0����,�6m���Ib� ��JK�yUh^��9���E`���K�
��Q/��V��T�"���-� �Tn��N������Kl��t�_G u�g����ŋ�	�!���!��>N@{���(���/͡�CT{�O��8`J� gڜ�N�ˇ"Y�j-ȻR;�\]4�ᖳ��կ�B �O�������x�9-G��*Q��)g?B���������%� ���L^�F�ekY���R�V�������Fw��P!֌�%06�B�(hE����B��䣆H>!���P����"j�����k�A����<�Q�T���IMk����N����ό���*D�"�v+�d�Wq�_%�.ƇW��|G�%�0۰h�x��9ڵJ%�5�B��W��M�,��I�j����Kr�A1g�L���N��ʨ{�8)���800qAʊ�]2�=�eEς�\�]>Dw�L��<M'CyeA�j�N7�����r��i��K�X� �e��E?lŌ���(K��gnȁ���Ϣ���!�F�e�%#��F�8�!����+㰓��#}H$��.��� �Œ��x�A�&���+`��Q�(3\�7�ɻpj�>c�d��sY]����[gL�+���O�,0�p�$��C��ҥ:�������dj<Zr>a��ɓy2m�]�΁-�@Jv�]�Tp��6l\�E��{7y����Y��Ն�]4�ʤv=���{v7V%�9���-�G�Z~��WkI����I�K?�#Y�(W�"���#E�W3��(����y_�Q��s�SJل��E�iOf��+���Vq����a�?i����qk���L��5
�]'���G�m�n��_�9�ϟ?���������q�a��_d���E���#�dv�B�����ctQN�jU|Gb�R����d�q���l��%x�{"����*a(h��ؚ��:�g,9rŨ���.�^��`�'���s;��A�B{�Aϔ�DfȎh���V��AVk�q�D7L˴~���Er��Ǭ#3���4l̓(2��k���:ήd��c��DI�7��|�+��+�V�o��f���`�_*Z|��5#=a��*9{�"UxĸM`^h�"�s%q>t��?@9�i�t������h�rfgM�	i��kvNR����Â��y�Y��z�_��c ���1 ��'�R9"�>�Մ�Dq��� �&=~�)L]Dȼ�BU�Ca��b,�}��R �W&xӆ�1+zh��/���B-C_����qtبMs�t�b��-:�w[A,���w�G�[0�f��s:�+�O�a�u$�j�bA�d���c-�A�䮉*/]����R�2������Z�f+r)WI���V���*'����� ����+}&W?��#/m�H+�aǊDt��=���}fcڭki�m�eR=�P�]��0�%��Dwa����X�`�`���\�*د��@�,�TڜT*y��8��vR��Dތ��vky I1?��ۍ�Z�Z���	�=���9�,��o��#Bg�s6`����`��(gJ�=��^/bƘU��@_j��\.0�au�D�W-/�.܀��W~�RXΘ�\9���*�B�a��?�ɉ�H�������}�\���1F���׋�+��I��8g��&���������GZ�7uLۨ�Y�I�G�d5Tց��.�d����,^cl9P�5������Ҵ���.��n���T�̓��+"[��lAܣ�3���H�� ���!�UfBّG��K`/�Wc�P���!�"��ϔ��X��	�i�\��2/=E�,�m�E�����APR��$)�S��<��LzC�ؕ��/�Lϸ�����z� O$H�������1�J��7�Vz���c���
�b�9w�IC��[��#���{��t���e��+��$4�mO��Q�����i��ܶ5�6�P��4���T��9��ehK�����A�!Nt���*>y�:������&���So[x���lz�Ko��B�������"v���)3����Y�$Zy�x���&+A�"��1����
bh����Bx&@A��B��:���g���澒 �i���<�����`�^$��?���m���0�����߫+>x:��x:�Mf��LMWC�(G}�*�\�;BE��Z����j��,��WF�i�׵��cE�y�ž`X4S>@F�-�]�c+1AE}��Ks�Cm?{��i�}bc�@�%]X��dÄ�Y�i���rS��Ks?����:�j^l�BlzЮ�t�@XTT_?.� 9��b�����1��O��`�U^f\�@2&��~q�&ҋ'��勑$���:a�Y���H���W��lB��6�``,;��v�Kn5yx��e;���IC��_Ԩ��:����6�NFXz��n��̱�z5bn���Q���@9P�3�o}��B)���>܈ʫ�]ӂl���:��3�lk`�'�v�-Y�Ѵ���� zv��s����f-����q���"��I�ʀ�[#�>3 E<�wc*w�-�>�����䨱�h��^V�=�s�K+�.@˝���+����$���f�����f��7/���epN5n.��5`�۹�@^g��%(��=9��of`(qo�b����ݞ*�xsc��Z��q�{�8����d��-!����l��S��Mp0��Ur��Đwy����m�,w�I�F��&�������M���h�d�-�ZL�M����pɥg�RW� �v}���&@�wOb9�~���c�7-�ڟ3I��f�+��HF�h-Ӯ�K��,En`��GI��ЈN8��^�/��I�E���-�1W9dgЕB��R
��~����d��4��#]@>�Ǎ�>)��;�`1<��#��0�ha���&���j�Ԭ�'��vsJ��U�$$�-#��=mP�ƛ]UT�����C�@&����P��d�>it
�"b7u�����!f9�"ө��(IAXch��f'9W݊�/8���Ϫoﷇ�d�Fq9&4:a9�,J��XS�y�녕��O�Ғ��)Wɰ�b4�Ԣƕ�˦��"�>�_$��Ї���i�_~������lҜ�c�܄� Sa�ʑ��Y�Lמ1����GB�g[������r���U"i��0��)h�`��\ɷe�JG(�-0�|�e���$��@��X�X���f����~y��%�t�wu5��ޔ�-N�O��!���"���q�|�ժq�~�{�֗��!�2L(�xtU�2>d�N�T��E�gS[m�Φ4��͂hCm6N)h?+$/�F���ao��r��׈2!�8S�z) 1U��[���%������G�xȪ������t3�B��.}�	et��`���-�9����X�����bt�e�I%]y�!�U}��|@r�P��*ezj������z�6!�{'{�T�H՛3�<�U�2��}f�W̋�T�2�r0V��'�7�mI��E���*�l���oɀ�m��7�N]H��[�Ъ��T��MjE;��O������'�w0l,O>�!��E6������*}�'�Re�o�^���'B�����7���/Zz�.@[��l��b�oPٜ+� ����!��<�t�-L��γW[O�q�����hp�0��$aT�7gC��,�a�8&=�ο��?Ʉ���^��t=���@��Z�\�~I�#u�E��wD<�����v�rʔ�N�824DTE�u������Hd=��m[1X�0�����[����M��!���O~ߞVdB�=hI*Q�'⇐�N��(Z۽;*��$X���3W���f�ӄo2{�rQq�o~�9��ZXdNPz�������,��d��)2�ZA�`�1|S��ga�#|����e}:���1oX��/����'H�9ǝ� h4�Ġ��&�'L���P�C\��l����
�H>Ou<� �b�^���(�Z����u��8�T�R<&�i�R�Kc�{�3���Lx�S�nk��:F��ri+M�G�sV�ߧ����V���!��#�
R�?��k�Mg�9�X
d��߶R����2Oh]R�E����eZž����S��	��PҊ^�Y����{"B���D�`wR3���t&��%��}�`\��D[�`��>�p��A8�A�#�*c ��W2���`�v��]_E�ѝ�6�mxz���yR,j�
���*�e�/���Ս�̔�ơ����Ϋ�()�h��x�Ft&8�0~x�����j)�g0g�?/��������u��~�t�a����5OL�GQg!c�[��Gm>�OO*D�������3�|�|��'0Đ��'b���`�-м��;/��워<�$�:�,b�7�I�X>�ʖOåv��	�.�6A#�,�2z�[�R��-�R�_��,�z>D��[�rty�!&��0�y�LHeU��Z*��5����k[���5�O�S$֒�bx�ͼ.v��v59o����S�%��'E���rU7Sq�]Bud��9���[�3�����`�&Ԋ���<N�� SN/l|y�7����E���kBe/_���bs�u��Ư�H����%T%��i�Y�v�c˅f��E?�}��R_2�����6u�M�G?���$*Td�f���ɓ�UAVQ��/>}�78�/�fUkMPr�l�<AM3~ԛlHR<4���12�U�g%�{-�Bn���ϒ6���c��A����#	�[����K=�������	�#���;��~��V1r���sӳKzfo���2MwM%l��5��P>Q�LS�D�u�p���}w��f�O�s65�}�����f�m9���	1(���з���m9�)�:�X>g�H�3����R��:�?��i�\Q�����l�^� ��a"(���S�:W�)�#1����r��,��0���d�	HA����\X}�X����_�{���Y3��[���D����LԎ)AɎ��FQ�%	�u��޴��P�5�����s+I9��n�Ͼ\y��2Y�+7�i{t�����p/���>��;a�5�"ӫ"��+E(ͯP}�M�J\$��� ��A���Yq�!�0���3�Q�aS��4�X���:hY:~�����N��}8�//����=7$������U���ۼ�0f\%��#+�مl&E�g}<�Ii�bJ��.?K�LL��/�dē0�kG,U[TζƇb��E�������m�.�Ӯ��H@*�İ��t��S��bG�mn���y~5��#��c�F�����Z��X�E�j/R+B����s�jy�2ԓ� EQ�۠��2�B�&�% d����P����j9F��|4�t3�b���~@[��|�N ���m����޹���3�щ�an�Yz̈�MZ�`@����Be�	�'��\%L�,DAd�YA �9�i��Z���υ��L?��a���J��`9�5�i���1>s��9�����٧|qZ&�d	*�wK-�<[�8N���F��ݏ�LP�Tŝ��W�7+��9F1M<t�i��N&���	q��so�x3�8o=���g��V#�����7l�������5&��%I=8�0�&��PQ'_ ��n�E���#PV^ 9��s����Fɷ1;n������Pn�&�3s�@դ�!A�P���,�5DfD�\��Yi2��D�f6KR�C�G\RT}d�q���E��(������p�����MN��B6��b�Ԇ;���~�uLW�_9w2��M=�;am���l�����)X/�� ƍ�����z X���p}Oѱ��l������_#���ݩ�%g���D�M>�4�"�v����>'�!����w�q�^��T@k?ش�⁠ɖ'[���˞ug�D6��4�T�3oW�_G�p޼��e��^�Iol�ļ��rZ�#aL�M���i ��1�����ߜ�^ix�y���F^> �R�Z�j�����x@r�������fm��[�@寈Z�5�)�u������G	*O�ƨ��ͥ�6��W�pE�DE<4B�t��:�i�]�S�i�3HEnb���~Arע�nk�Z�i~��V�;8>X
��,���ߨ~;'��f�x�x��dU>�q�s�jO���F(��4����=Ld��B�6#�&�NH��0¡�̳o�LMB$�W}'Q�a/�|nv� _�d�����?%E�ӡ�
CD�9w�P��Z�@��|ߙrˢh�̤n��,�q@�22�P�ʉ�ސ#~������6.������9]�*��s��x4#�������)�*��T�FT"��Q��l�?ei����12z�k��]1�JldfQ�mp��>B�:���+ыY�Z�ޥ�[vW�Z',�~�e��Z��B!�3r�o2���cȐ*��`��ݛ1l��[�*�d��h�i���enj��ۡ�>5&Ԙ�`\���0��|{�`���ba��[z�S7�Z}����^ޤJ͐���0�(%��3�(�C/GK3+��O��Y�Ɍ����8���T׫r��Fdq6����?�cΔQ�.'% �9o.�0���C�ͦ�DR��Q��A ��]م���`��F/�OR�]˘秚WS7�\9*Em����=Ql���\���ouF���ˎ�,����ҋ������<��n�λ���FCBQ��O.Vv),WrZX�-�����B␢���pS�>K�]v�3���Tl�q��x�D����wq�9[)����l�+Ł�oiX�['���0-ns�ܪ�i�����9)�TN�5�~��qt�Wj���Y��C���jԝ�L������*`7"8���"3~9b�$��pU�.��TS鶜����U�U���9|����r�d��u�8e�H�P��RsU&
}���th�MYW�`�%N}���I2��:��VMIP$w�.���	t����7�[�Y��&S��GʺRg��c��c�`�(��4�+��
��+6�����!㸎�*�����!5~�ޕ豘�\��ğ��<�r^T+�b2�V"P�޽�gI�n-5�=��Qǲꛎ����/�e�A�����xp��YH����Q�	���Q���k�����~��c#T��'�7��.����ִbc1c�|���_	AYL��dv/��U5�DJ���ݞq�3��q�Z��Y�P&�w%
z�2`����wK=1΂��<�A�tǒu�^
��cf�r'{9ոƁN �R���z��E:b)�=m�SyǢ�.���56�j��U�o��'J+�0r�pvq9���u���X�F�=Y��H�:ve����qm�ޜ�	*�kJ���(@u���B���Z��A%��Fh@O{�^���Գj$�	��`'?Mi��AcDG�pQ_x�0w�������i{ z6�ৠ��W!�1X��U��v�W��������߇Z^\�͂�$�f�wia�jK%�?|����l�#��fQ�pg�F#Xqi���	�ɉ�<�n���8��4ү���*���7�����s��&�M�"�b�Aɭ5�S�b�M��	��Ow�o����
��G�$�ى�7Q3�:�Ua��ӕ�n��S��Z��M��u����̵��cE�K*	�o���j�cS����1�@*���^{٬V.���3��G}ƫ.B{Fxٓ�q-��Y7�] � JNgұ��/�HU��VS��aF���`9@{^��N����*��������=uTH�b/j_�f-ܬ��I�������>�,��|�^1�hb_	7���(�k�Y���^�uo�7#b��q�Nt� �g��1�管��~p������w�4��S��Ţz'�<�!:A��<�#��p�0��/OU�?�������\�U�#�u�+{��XF��K �nm�q��m��A��H�n��{[E�[��^���?�J�`�d@P��f0�(�0[ڇ��9���q���x���u1w���U_��x1�'��U�{� wIC�}Z�T���&`��D��<�̙l�Lݿ��$�1�M�����c�w&�[�bW�����_g!����`ɀ=jمH����m�m�(_?;>�=ޥ�ME8�R�xYl�^�L�V���+�j#{M�Ĺ6@԰������V#�~F�Y��Z�J�C7��m��n��U�{�Lp�y^2���[d�u��^�^7nd{a=���	#O��^�U��}�j�Ǜ�a+�J��6#����:AD�rS�ê���׌��S� $sQ:�C�K�S�0f
�<~D���맄����~�ۻ�1��|yH�������60��6ok��g�d?h�;�(���S3FZ�4����cS��&D��C��%���H �01PPAx�,�?��Ro��#[�@O�3����Z�Hn��y��V� -����Ok����`�f���j���d��b�-��Ǉj	�K%�o�C�2�Z�ԣ��!ĺ
�u�f�����䃉eY�{ #��ϕ���o(u.��"��R�h
7���0Qx��2V��lEkV=��r�	�9��W���@�0�Z��xQ ̅HC�&����$;d�F{)淤e1r��	T�Rae0\]��ǜD�Ζ���`'�_�*i��Uٶ�ƻ���ɪ�Ͻ��]�u-�3�Vј_�<&g�`^�`MDΛ��;�ˢ��	AέC͎�޹kE�f��s���٥�D�'
ÖZ�~	��Z��=��xt._K�_|h��'��]Hj��8�00��d?},���C��F�E��B����挗5��X���Y"+w�85���ԃ��Gs�\e�����^J4]<�+
�t{�w��ȧC�+�`NŅ�#�B7p(�17_�����r%�e�N��l���&�볞�e��Jm/1��&�A��j�����#s��A�3kt�|�z΀���t�^3���J�'K�%��f����%����˼Fi�/�����I�MՏUs����(��X=Mu
RKN��� ��׊���O4���\\����r��"ׁ���_���}6��wl?lh ��nWpҌ�uCt{�4���-�� �>�%�6��{�2X�$��^���n�4߾W2V�o�۩�z&5A��n�@?,E.(d�A����|��=s/vl���2���T��/s8�ODW���w<Y��3O�B����O��,��:�Yʃ�B_u?<�E<�����@���ni��h٠�-ɾ0����l�F�,�G��u��o��!�ش9�
h�@h�i��U�n錎��~������	���N��c��Xa6���ঠωXlʖ�߀���xA�gX�(A(��L���66ԍ.-��ԻP�;�Ty{��`��_���6��u)Y^��'��%QJ �����Q������M4Y�/T�t	O�4��4A��ð@k��n��:��}���|d������i<o��
4�:��H���&r����6^���&wo�[�r��|�0I(�˚յ�+Qe�IO;z�FZ�X�9���儨(E9�.�a�t��?�%�@-�f	�i���4U��o��r�X��P�>����6gz�t�{����rsC^��@��Vڶ�����^M�9�qq�ӓN���m:���vv�B�����;|�b�Li��Q)�g�.OX���290���ԟ��K��q�X��뷥F�����2�0��\��\&a�³4�.���ue� up�m[V~���I�'����Z���"ATJ�HH�O{�S���6��	��Z`��l��k4ɳ����R��f����3x�|��������l����9^'�#���Q���+�ed*�շ�����3�;W�.�*�)7��E\)��%���Q�r��is_A.X����c?�ʡ��s�z�Xd6���u|�eb�)���ە9���`%��[�u><(��`���.��"\J� *T6�� r	�������8�����ʜ]���h�,{��&�]��� ���R
*B�bN͒���~��K��:wEz�z.�a�?��,3����	�`8�N�(���k���z�*Я���z�fɹ@�$]�"���`���e�E�ݍ��/ ���5H���v|ϊ��=��o����l��5��zl`��%��m"�X�G��1�l�;�׏��Q��҄cU
L��d+1&�����}��$D˺AWE�W=��Z�$��+��m @�{:�O��ׇ��Ϸ%�	�n[	���T�Os��]�`V��GQ�j�iI�|���y;���7K�7���p6�-�C�F�\W�;L�hv3w/�Q�w�'TCv�M��LD���|I�E�y}tR�}*���0���	���<�H�`�_���t�C�ڦx�d�N�I�Yf��)T��Ig��;;R�ch��CzJJl�󐜖I��c��d'-$T�ڌ[�*J��G�䱛
�;(}Hل�l�:�wR�n<�#�@<��q=�x�!�e��h[B̭�d�>xǵ����7��ȲӚ��x_���<��Q� -�N�����j*�!'���ߣ�L�ԁ]�������8\]�� h�]��ۆ��EK�� n��?�j<ƈt�v�l�ʉ-<o��^\)�3���n6�/^ ����֙m-\�`�s�:iÅ=��� ��<�o��E�|k}[^v�O��땑3W�Ve�'C`�֝�fh���H+*��;@�2�;��-AA10u7en��QH��\�B[�|lw?U��Z���CBzt��I �R�! h:n��	vc��Y9�����.(��K^�eA-�t$W�1�^65�6z"X���q��HH��5�u�$��Bo��$�?)`�Ű�jp���Cܝ4�@p�(�p��+�!��Wܻ���E=A�
2�A�����?K��Яk���Q���1�I|?$-7#5�Ϣ��L �/����B�ٷ�=&
뽹z�x��j�f+���n���0!P���%Ӱ�2ف������u/c1�#D�s��*z���ǘ �sy��YuY��u��b�so��H����l۰Ry	A�[���Dt�b����h���y��/i�{�k2��8ft�fr�chS����,N=	a(w�:�a�����[K_I�_dm�tF�r��`lf�(�ՃF�A,��=�r���3�)B�}W�3ڋ��{�ʝ���5ϧN:X4�-�`�Q#���i�h+r$��H� V
T��*���mаfK
&h��7�"t����K
r�&�d�80����$���r%}��A��U#/A�2��cE��*�����^?�u�LZ����d<�8��4�Q��u��'��C	���<2��L�앫+RFs��屿�����I��G|\�G�f�醭
I�$��~C�v�G��h ��]'$�q�{_��&|,v����iS��na%i�&�]
���n%���{d^b����S��R����
�����uI�zaī�}��55C�PW.&Ӗ���ڇ�ʼ��͋P�Fn����<4x,G�e�4��r�e /wP��A���WB�A�"W�5�x�;��'kt���~��
X#2p�y|�+���~4&=�����V��y�����E�ۖm)Bu���i2�FsIg�[`��|�T�@����9�챏zrʍ�+9�L>���?#�M�a�k���k.ў��Ī��?�
��;n�Tƪe5(��F��vx�"{���0K����Z/�B'�I�����MRW`4�baɑ�B��
Q�B6�Qv��Ȧ;�S��ah"�6��avB@,��
[e���2�TS�k9�(�B�>�#	W��sk��
+h��P\����a���uA���o-c�2R�*��%"�-�������t4
�S��АF��s�;2渪�������g���v���Ќ���es���?�PP�?�F6�Ҡ�B�K��O5W���]>��K&J�(����|�L�i�xh;�6�Y���U�dT�O>����CBӏ�pT���U��šJ.z��i;>�4h�1�t��ʴ����t\XZ�IZ���=+�xs�mRy�8,R�(�E��#�����r�:Y��$A�>}^�z�N`O������&xS�%Ykh���*��B��+��9y�4���[�|�f��,W�3C��J���H£`
�A�H�Y�����{��
��.m�/`��G��"j�s�C@PX�US*��a�8���A$]���b�&D`���=���:��ւ=qP��o�'Im��F�fl�&��c�'�\�	�	���7<�y��)�Ғ�J��>���{)��f���BL�@z�i�I���C�@��
o���	�P&�?�	F�zqz�@?���i@3���L�̅�5�|�Ak)�nw�[-D؟��5��Z�W@�誟�	�W�LO"oΣ�t�cЛ��p�_�ǁ��1�ޮ���EFN~�����Y�YZ�KJH����[�/����Ћ���u�7�����4��rI��Oր�:Y�C����4�h�5��oU�8U��#�:�^C��t�s� L&���:L$o��=�A噩�Q�d:A)�[��C�T�i~C�<hP����FF�%xm���O�%� b26�hKk	����=���N�VW��H;g��n�c�H�')Pr{5@$/�Ӭ�,6�XI�D�O�v�<6�d0��� j��Eߑ���Yx�q�ҷ�93�	�Ŭ2:��/U���uU����%�0�L�3�h��	��Y_��,t�~LGs�-Ǽa_u���榋tPS��7"t�f1�RX���p;��=�D����U5G3v.�`°.z�1W}hya�_m��0~p�`��IXLO�����Ѽ�5�/��)����5 �	R��*���'x%^k1�T�"|OɈ�J�|�U�Q��@/�C	�Zj��*�}�'g�>��E^�&�H�֬a�9��W.��x	���� 2�>��W>Vpu|�*��cd�+1g:vY�K�����T�Η1��R�@���e�on��q<����C�G��eXd[*$4�j)�hiQ�a��hR�	C��OWHʈ,L�Ԇ6���������L�,iSE��C�A�pb�&�;p��(����T	��Y��q�L�F���h i�ߴ����9�@�^�t[&�t�ւ߮�'/�-��|X��FI^b��.p���~�dN�E��V�ƕulY��(�G����������:7�<���uy�-���Z���D�Ē�
�.��%��,������.Ȑa��9�A�"=�o	�^W�6ߦ_.�$�|
U��Go�?=tK@�S�q�+D�݈�@a�0)���rE��-�^`v�hm�c�����;�ZV��Kۿ�x�����uWr�iت���R�q�8����"`���Hmfdӎ��0y�^�RB��M�Ƒ�����<S)pj�����ǡ�������E7�?�S���3�(�X�Z�͚**��7Tx���脮����*)�|+��L������Uh����b�B�}~ d���n��Z;�>��Q�0��=H��x�K�){���_�5��� WxC/�֖��q(Y��a����?�|����ߤe9�E���NT�����c�I]��c�0��z�A��|�]�D���R�ԔX�͵?���/���}���AO�ڛ���az�������U�Z���@�^�0�[RK?($�_�O���]����J�~�a�/�����s��x�o�te�<6�Y�}#^�>����Qr~PG�=?�;P�2�����8A�y��+��*���=wdI�
�:�n�=j����|�ߋ��?Ev�[�C
�^���ʉ��+x@d
V��)4qx�&�I�. Rj�D����j� <�}�\6�DM�f�l*>�!�A������89�v1tiHy����Q�ﴵQh��>܆M �j���y]z�GW
�_��!)l��&㚅��<�֩1�]E��ڄ�'�wU�C e���AG��ɬ}��`2S�T�����c�����	�a������JcH�E{+F��g����d�jO]�H�����`ƒ���䉴�ڽ{D�gF?@v�<���Բ󾱠�^��GT�F+�I������p�1z4;�ͫ�0c��Y����)��.�茯m/�s\l�쾉	�������A#�i�8�+"]z����#R._��),��?�-�a�����+Q��vJD�d[`w'z�>s���#
�_ҥu6��~�f�	j�����`eU��n�~�;�R'�o�8��\�+3������
>u����+���PHS��pK���	@Ȇ��2�W�'��K�mڅa¹�o�U=kk��qv��`�|U��#���]t�bgEZ�_���9��	�l#����V��;����U7�&�3dq,�L�,DyZ?�g���jFD�183(|�XM~M�y�m�M:TF�m �o��N��ҐQ�b��5^*�����X���F��C� ��d_!oI.���
V�h�;?!�y����ޫ6� �ܾ�����c�v>Aĭ�U�^Q�_���)���&ϋc��Y	>2�S�0�:ux����H4X�I�|�N�^R>^H�c�J.R��^��v��8#�P�m̐�Iн�qŀm1�-���'�Ҹk��� ��H�{���A���%|��I� W���x�{�<b<t�	U�N��|=8���V�g��U-O�t�3Г2��sLn�$��+����<"�<|�ց��*�X1���6y��԰��w��נM�vY�_x%�h�7�$T��E�%N�Rr!#�%��[1�*��(˱J���ǒ�:����z5>S軚:R��r↠�L+I?Ã+�ݯ��I������W1ݒl�W`�F��@FC��i �,�I���^SL��DҎ���pϢ�E>�U䂙�|��5�x��y����Ak_��]V��Pܼ)��kE	L���M뒏!��K���^�:EUE�B������|���ٰ4�gުd����� A
�������Si��.�ơ��]���d���h��3m��Hv4������a�g������g����%�%u�"�B�"�T�s��q�o+3���X�f
�U:�G��u`�:hqH\�s�h���;*x�4,n��B���=��mAX���f�^�z�sxũ�4�p��Q-�\|�zt�{h��m[]�E�5nX��u".���'�kJ��1C��9\ti)'�iԕ��5�5����sdH�G4I:��配�yŅ�}�� �
�Ep��U���ٳ�4B}��h���������G�j�
 �U ��UB>�q�����,��_��.A%��nbF�2�P6�Ϙ�!����t���	D���M\n!��5�ח�r�!N~��8J��_\��h8�f�Q�O2����܄�8)p|���q�<)Ƚ*»7�p<���¿�@�����@�fjZ�\��<�\��)`*�Ǽ��=����Ѻe(l��<���l�����B�#�J/���2�Eu�p)��ݙƿ�)g��gZ�{�SI������!k�����&���S��&+K����`���R��9���O��B��m�6'�������jV�En� d	�
���H4�Q�ہִ��.
��y/����B�J�2��R�h|�����(�R��$:���HM�+�r� �M!�pq�΃T��+D{~u��ښ�9*��ZយE�bļX@��`f�8[�C&�9t�%�)��>}]^84}�����伥(���:��N�Uww5�!(������;���s=YG��Ioz����}ON{?�����Km����'��0��<>�5��y>[^����'��2�Ďh�%
�c��K���^����r��S��N����XU�.�Q�ۭ6㸤�k�苩���cJ���V��Uxn���x+�M������1� ���x����`��N����)	���\�ӱ#g-�lq'C���e8m%��b�g���9��s�%{��l��Z�QB�t3���n��<\������[BK��;����$run�^nu׾֯�y��(��� �2q�Ga����ko]��
��<*N��67EW�o�Ud�?(V<e-��O�s � �(�,Ֆ�l�,{�����+��� )���U�l����U��ɖ�������`AR?OG�0�׷K��1�I�9�}zC�P�ۍpRy��jm,�}� �*���P<C�=1��f�� �{�+��K�P't/�n��R*��LuЌ��Q�J�-��]X��}x\���܇��^��F���%�5�b�<�csn�0Rs?/v󉦫�/��	e���3���Oh����M�4�<���dz`G�CӐ�<���W%@MJ�,���ܛ���ꃖ��4j��]��ו�fǹ�D����Z܉x� �{j� ��29�m�nܚg& �V}ȕCA��J���ح0�8g��;oϪ��i��~ U�|Dc��R"Ȍ��+�6 Њ2�"�XU���Y�C�7|6s�K]~g/VQ���]��O� O���j1Co���Č��A���>�	�K:ֺ�l���@�ZI9G}h�� ���G�..v %M+f<9��������7�b�*��NV����`��}�<���7@5�lE�"L�u�M�s�Ŀ�Kk����7Rm� l�ΧvX�B��n��_�U$ �D����ӫ��G&D[�A�����4Jxmj6�S[<q??<NA�����[�����D�eX`�qa|��h�;�g���.G����u*g�*֕��]GB&�[�� �����:���>K���ј�S�P9��>���0?��8�}��f� �z��F�N�6���LH`k��Vf��{\�Ӏ7+~IW��46�E7�k�o*;F"�]�%��{�6Ŋ��4�z@,�F�栬nK�CAyQ	�pش��3�g��s4Pܑ�7Oq],�����T$cn����<)����f����V\!}�{�`��t�m�i^�x�s�����=����<�9�s��ǫ�= KQx�h%����݈I@_�$ 2�@����ʰ8k���@K��>��=7�5K�֐����
h.�I�=��Ov�ڗ����J�jɨd�J�l��zl!h��&L{�?9���p��ְT1T�$���$�K�K��	���>I��L�$2�&ʠ	��9�� �^k��/[�H8v�yAˑ�g�x`�O�ŀ�c�lFN��Z�E*�3냵�~�t�w����Р�6W7��{��lL��� [���}��u0!Ln����t+�56��v�E�`��&�F����>��W�D������Q�*/��B�F��K"�r[�J�2���ST��ԉ��)�Yx�Q�[��]�c���lOF�E�V$	@�nO��أ�}ȉN�5��+|v�܆s�s�<s"F:A^�#'0���s��"�/�����Iu�~7妨��Kl��,5#��K�7�%�xY�����$�-�+��g%��b���#������{p0��4j*���lӃK�����D��侀s#~��bF�	i����i����S�d�Pu��b�%�f����Hl��U�Ĕ����Z�Oto�<��6W� ,f��������L|��#T�C�R��ڽ'ܥ�r r��7D���L5�k�B;d�'^�6�(i1mKP��o��Z�w�A��|R {���OEcgt)1���c����[~�m�H�l;S��CV���}����#��!�45��:�>M�j�vo�1s,kc��@>�(؜$���Zw��N�&�*[�g���y.���]�`@ƕo��'Q3濏�ddȰ,A�����C*�x+I�G��>�6h�Y��F�7 �s�y�msV�DQ�~rW�A!Q{,Y�R��������Y��>�ܳȿVH�~���ӛ
��3���njU{�*�Ly�⟭Y,~�tq�$����f���3�/�פ�	����h&�L~i��@A�#H�?���Q��唻�#Ŵw���qE����m��>���(6�L��"�ƈ2&����J����&>�6��INfh����b��h��k 3�Ah�p��×�~#��*�+;�?k��=������E(���lVa/H2	P3���Y.At(.�~%f�B��}��X�I5��82ϩ6EV�eS�:4q�� z��`	���I��@2����k�lÞ�#4��oCͺ�TR����.YB�J?e�k��L�&��I(PO`���x�F|�¹� �_fpYH�ؤI&q�QN��o9=`��[B>���Ա���jK��ZŢ�ۥ��E�~��|Po�=&{��ӺY���\z�MDh4���Z���y�I7�y=E����7@~��&|�Q��υ��� ��I�{֤�oX���6.����]̳?��+w�\�bE~��%�L�f�."�9��~4��E�D�wTbxd{�|������uo�/�� ,���D�E�&7y>=���6��\dsL;��:AŸ�c�����fP�7��)ȴXy�W������]�k}�C�8�P�r�lz��d���OJM��GscgHb
��w�$��?@�Fr\��3����>����8�������~4B(��~ݻn�P����)/�JS�����%�9t�2���ZpO�о��դ��?b-������k?�@�����N?�x�/2��_��}���7� #��oo�꨽��D�ڮ�X�Hm�����ْ p< *��X�����yҌH+x�5�!%gq�L�AY�XY���
pD�����ٛL��Iৱt�'�����������$S#;}���_�@.ݭ=~��iL J���z��D���l�o���K'�����:G��1y�����ç m�'G�93�T4���d�yp)ώ��~����Q[��9@IH�z���s��
#�)�h��>�T0�M� �������-��Ȉ3�<��h���ͦ�ɉ���	*�[�G� jKI��%,B7g�GȺr�A����nmD�%�dɳH�3��$CK֗a���3���X��_Y���y���Lҿ���qЫ�KNk@{So�y	��unMI3�CMi�w��w]�l���9�IL��zp�����S�M����L��sv7�^��*y�e_.����/��_X�/G��乂���o��h����Y���HR|�[���T߆X�,;6�����k�6�Ƹ�b4'�^Q���"/zh�ի�CyN���pg�$_�n��l8fAoi���E�5���P.n3`�:��je�~G��ӽ�4�w�N|��o�; zf3f�SL��{t]3�|���:����>�*��ޣ�xh^����?z���2�E�;Cӱ^bkA���W����e�E����r ��9Q�F�'Ĩ7E(����yv�G���?�4�g��%?��eM����WNS��E@{KA�X98�pѻ�N'?�	�q��zޫ�>�Gs��޵nU�*{>)�(��?���f����{�p�M{�}���һ�HˏΜ�����$��T��.�.�"����&Jd2���U�$���3��>���WB��eԑ��M	6�S#vMYL2��0���Ћ�r� Qi_��ӡQ���$}�1:I�yQ�f�.�]ԙ��-�Vȗ[�e/�J�	/ɜIUJ�3�8�J��_@������%[����籭Z�^�~bVH lV��:�Tmad��4�1o�_����׿� �B�HI�l@0.m�e� ��Ĝg�:�{�j���m����G>�.KY	7�}:��`�
~jfײ��@�MkO��52�U��#�Y��|�^���"�w�� ,J7(��uLiG��~no�	��s*��t�ɶ��D+�Y^+M"��`��R�%q�On��M�|�����]"�MBն(�=B�J�B3k�����½���i��h����޽}N�s�A��$}���nL��`�{���ZE��7�l���Cʑ �rg�Q�r2�U�gĸ�p���Q�b�}Zo�~i�JQ�^y�F���Ck��qi�+�_&Ђ�8�tΧ���.o�YB��S���m�bI�t{���I����'y��&�7��= Ě�ZJ�c�G{�R\��:E� ����k(5,��	���BX�����Z�≯��a�6:�JEY�Q�t~��)DZ��.P��!b4���y9�l;cg7�ǡ���caZO	���* ��X�	ˊH̎�l]�[-gU��G�Z�[&+O6~O�q�f+����L�{a�&�O��Ą9[��QH��@LM��p~��	�G�G�����1�+�a�2x�/�t���0�֠���𲞒N��˟!\��C�o�Y��pK~<+�V��j�����8�����5�s\&ב�S��9-<�GO���Ɇ���}�*aB���5��{�A���zw�]#��¹\�L ���1�$f�ح�ba2��v]f
�=�����_
�H��$'Q��������4��)����1���ɱvm2����B	[zv���~n�T�Pώ�o�}���R�ʆW�0i�,.�iJ?+d�ժ�N�?I�^m���K���ڏG/>����BH-��'Yoz�-'�zm>�#e;�g@�+�`|�v����(O9�y��w�b6ב��N�R�͎Y��c%%�y/=��%�^��V\�ZeJ��|1_M-Y-�� ��(�4���Mߎx �nK`fx�%��@�h���wI��h�q�0 ?W�;Ŝ{d��{~7�Fhs{���Z�4�ܤesEm�^�|�����1v`~`�ڃn��%OM��n�޸�
��i�X�EL�d펮�䔽���t���i��>s��+�rq���-�^�a���ۃ��c ����V�B��PV���V����Ե�?�+�����"n�/�>�� �<�6���^z��'�"L��J�/;\Њ�����s�
� �������X	�%��K���z�p�xQ��������`�Ku	��:��ȰHw�ŏ�o�:9��Z�$����Ai����I�n
)�A���ķ�g��`՜�c�Dp���AM�=rê�T������������w����	Q+�a瞠���W9O�S�Y��/��!�Ƀ�i�E2�0��|�2L��<N�k�HX\������n�9N�2�����!!N���b�� =�{\����R�8PR�@E��G\��!��H��UQ6"�iX;�4H���Y�>	wxp�x��I��[�������G���Noئ Lr��@���8��(������_�e[�Nn�A�hS�O��>��aQ�E־r�Mv�
k�+y�q��K�D���]=eK�ݴ�9����Tϳ;�ʰL��	�����6±V��0��rk�0`OQ�k`ƖI���Apۀ���$�^�Wa������F��כ��GVX�'�1�TwQ��<X0��c�ZS+&�P`�T/�$�OT��Z^�q	��K_�Y�����ܗ�TΑ}iS���Ê]��p�x�3Z^YA�դ���jQ���j�T�^]�c�36�t�6I����>�;�i��������#�ޏB�k����-k$W����{�ss⣙r^���/�]�a��N���*�7t~�I��8�'3������E�Bs}��qTr�0�y�pֽ����ſ��I�l���͸���@�1�B.{���Yt����t�s!7)�s�PPS��\%���'�,e���w�ѥ|�X r��l2��<h��ʤ�	Uf!Z~}l���>�CH�xc}�b��L�jġV�Cxu,Cf̿���b0�P1�?:�U���Ap&��_G���e/2u�M�ӷ�d�E;��4|���uL/��x�!���0?�<!q�W��.�\,�S���e-�K��m�P/�"�?" �q�Dq6���QR��yJ���=��8������"��OY�`�%�ҼP�97���2]m��`���D��C�
���v[LwfD#�V�e=kne\;]��=���XB�ߔ?���7$&�o����"HӼx���]]gm({�s�	�h�X��֦@��1�*��.�6��'�ۅ�2��Srr�E<�[���CC�B�7���Z@�^P>: ���B�{����%�kc��q+��IB/�P4�*�̇h7�n�+���K~�w�y5��d6R{�dM�u��<pU�	��Φ�XG~^�e�����B�v�9�&T�\��B9�+D�*�F<�9��N(��~w��{� ��HOc�+i��6����9���(�}��@���Nv�&��C �Mei���t'�}���
����#��y��y��A���TW-C6�$� S �1ȳNi�}S}��1a�Ը��%�]]W0]��5�6HU�+O�Rʿ�Ai���r�s��s!�5����r~�H*<c�$E��¹���#���u
�7)��DRj����xI����1���U=|�McT4��|��v�T(	�3`��a�sfƺ���a%�'־�4���S��f�}���5��)�U�Q�Q�(�P�1m4��И�����;i8$r��$���dCԦ9T��C�%쓛_����R��<�\��v�F2&��-M����V��u?�ٷ�������n�a�N������4��F\�w�r��g�����B{3W4{%)��y���ҽ��r���or��L nzϿI�zR�Ԑ�Y�lMν�6h�*��0&)9]��ˣ$�Ymz���K-{*����:���}�����s�sV�]�����SP�K�~yS�i�lm��9E V>W>�d���8#Īx"Мnֹ��.���1����Fj����g
&Ϩ����4ۚ�+\[f�)�K�3�#ǣ��P*������8�	p���C7r�ʓ�d	�Bu2��������xڦȐDQ#q����: x�����3r�wY�y6��o�e���(��GS��*�ne���,��<Q���\������MgR��Cc�]���+�^�b|EI�5Dĥ�J�h2T�9���Y6��b㸋���3����|�f�)����fFL殁�l�+ƫ�Z}S7�,������t�~�:t��M�u�9G������˜ưD���e��d���ޜ�E
���6{�xY��넳 S6����@!�rV-�-�Ze��u����*���*�r�>GA.�� ۦ�����R]5�`&���4[R85c��`��S��"~���%��X�dϬ�?��y	��U��JL�ɳ ���;��TI����d���8���!KJM�S՝`V��QGxѧgI$w,�vML��ʀf=�r@<L��9	S�!v$%�ɺ^�s�{#ǽ��]{$V7��.ye?�a룠�;Mm.�`�:K?�b�R��O�VD��-��sy�H�Ȧ�I~%)o� C���)�B�=�� �_4���Zkh�Ktez�x�p��_`#�ǿ"��3�����,�9d�s-2�h$dN��7�@C��҇��z#<u��;��۔�y��5���P���~�*�2;d�Hl
���
���=�?Cݟ>��??�yg�h����wUnǁ���ȡe���?!�1���3���!�<���szYk����oo�=@*�	��:�^=wRYk����C3�]p$N�NLar��3�h��Kg/g<S�C��E���}T^��^�>�eq�^z'K
�������6'J��U�,��t�Ej���rAK�W���clp�r����ž|Ce��`7cٔ���~�H�u��\�lv���8�wǢ�[JQ���@"%ի8/H�8���H�_�$>�~s��T�?dr7�����kEe�5�gc�le�N1��M�����ko�0�l���
��yfp5xk��+�\�SG��(&�R.Ǌ���S���ܲ������M�=�]@�ޢ���2���0�	C�Ͷ�_QNV"��/��7�|���_�[i�=��Ω��bcJ�fQ� �ƒy�ٰh_m�C��J����"S��i�u�y*Mh
���=�L/��?�[*��k�/�5�?,q�ͧ���0�z�3P�)#�{�X�#*�i��W-�_�~�җN/\��#�a嬖U<��z��@���Yh,�t�����2��h���Q���_dq���>CcUj�����]�X1�Q~��ػ�R��a�0�-� 97��	�l6��n��T~�:g�R��E��7�z��x�t���@��w��]G�@���zLY�w��u���(Wzlt�ۋ��G��{@<��`�_�� ���˖oLk}�����V0(��\܆���Z'�{��P$�h�!�'�{k�D$]��/.�iq���ĩc/+4��:�Oǳ�������D@Ji+>��jņä�+�H�e��e2�����h=����H��a ��ѫ�\5�L���H��c�,e���Fp� ��)���W���ˉ���?��]c!�L[� Ӟ��`OV����J�����.�߁뫏0���O����[�ӢQ���B8�F��W,2�4S����-#ĝ�F�I8��q�w�T8m�^禒"C4
�ߓ���<�C�H�؆��\��<�?��-��9t̚�
q;����f*$���@�̞�}�>����A�����.��<����S��'� 6��|X��>`[���� [+��~��`M��`dg�oy�M����g���B�FV���G�¦����9��uF}����-�D�*U��hJ ��Pq{C���O�я�E(���l��=�Χ��/�R*g�C=��\�r�1hkT���:�)Q>�O7X�~
=aaH��q��e�����=N܆t��~�y�4Ut0"�!��^���&����&%�0�Q�`+2�@�fY��ϵo�k�`h�7�'�Un=���B]C��1���{��^�V�xfjh�W6�Eƙ�Ky��Y�Ey@�4��i�Auȣ���X�{�\��&  ����R��p�*���WL��y\��p�|�Ѱ�)����%!"�؁b(3�"��
�r�I��u�[o~E	����>V���ּ�Ry-�W�S��'�':�NԺ�+�SA���뫮8��s�������o�b�n��tg�v�2,�!${&� _�%��z^V�Ր�)��9�,�己���|����J/֘;�] ��m�� ��
^�k-���䖔iġڸ�)�X�������^�0�|v��Z�`�e��х�h�':�0�J�����͐�D�����7�g�A��'j�P�u¶���/i��W����S�??|1h��xO���]�ȁ����4D�ݥ���*Լ�O�c���Ԏ�*pV	�鉹{�D���;۪�}͎�3���C4Y�pXQ�����ҼQl�	{`�T����X�qە#��ȉ6�SAk�6�w���໪�7̨�/pԌ��ф�s�5*��k �x��r�L39p�8 �A�~��D�{y^W`g�ٴ�c0n�GЗ|e<p��y(3����{��r$C zCk'��@Io�BF.u�91h(�U/�ZBT��8���)��A
�l͓�%����GP���*~����Ϫ�"�C'�Uæ���Yf���^���z����3��}�0���86��3>l�FXCp���\�<[û�8h#�_J1�Ȏ�����@��6�8W/�bŁI�Ɲe�q���5	>�e�J]�ɘY8�8��.�e��]t�>�^ѝ�l�p�k6>7����2έ5*Ma�t��Ŭf�l�4H���Q��i�*�_+<���M�wG����O`�޳��6h	h����˲�80a�+�h�\���i���>�.��w�ꀷ�rg�j 6�W/u�t�l �j�"�6����X	Y3�:��f<=~�P�EC�
������Wd�l|�q��t,\��J�?���޹)���r����P��:�_��I��\��B��.'f �op��?��.s���Wu������!��s�����	� �:��ʩ܀�9�Y��`�Ά�D�cW�8$׸}���NS�M'�3+���hD�=�( �bV�.i��y]��G-��_y�ƞ��g��9�@�lӖޢN[-�-����uƎܤ�nX�w�l̞��+z�J����F�ps�؎�h� V�����$��nF�3�=7c��A_�oE{��2�
��)5�F��;�0�M������t�?QN#��91��9��S@,�)})3�'�c���>�Y���L@f9�m��os�BN�G����YL,�ݚd)ŎOe�p�?2;w�%�N�23�c��0�w����l���6��$�E��&����F|�uj�ݤ�0S#��~(`|��H1�C,��ڱM�	�^~�xG�'n˒V��!��l��=��9�$�KWv�n�ΡAc���׊��0&H�1��1���\̔,��'��XT7d�6J���FK��l��x1�'T�e�J+�zE��JnM�O�Ƞ��7URz�_]Kp&�_�����#i�-=-?��(�����zDí�[���P�pi����&��N�~�����^�5粽˔��4.4��Zj��O���0�E�6I�%�z����з؆�Omp&;��ڡ[R�U@!/�r,�dܓ��PMr��,��NkO�n��)i�_��DJ����K{Z��"�BbV)��s&{4EO��+F-p�R��g
0�F7qRH�����yNq8�1!�c�'�I�x5�j��Z�LB��^"i�-,Tc`�\�13BLv�͗�-�R���i#h5������P���;I��%i-��	K��yQ��x���f�8�`̫�����S���vi��H�[�U4�͹+I�73?���������òL�-B@��Y؋�����q�UY����+F0�"�ge�"[��Ki���:���<`�h%l6�)T4 $QG�>���a	�v���)��c4.~�}his7�A��[kE���N�}�&:ɧ<�8,�h?]�������e��4+|�B�da�E� څ<���J�\�Tp�}�/�6/ z������9�hٍ�ؕ�dBI6���w�#*d0�ZGAy��E���ZǙģ���L�ݠ���2�:����
�,��9�fV�+���s��t��	Rkps%��Zl��5g86��phT�y��+�V�nʨX������D�[��Gl3|x���iERj����@=�&�~�����?|��p��cO�s<ND��D]"�2X�P�SR��8�Rf�(��<1nM5��]�v�p��R_C������-O��2Jm��q�s)��c(�q�?��W��Y4�첡8��s�h�2Rf�+��C�v]�z�$P��k�d��]��a�MS��ѐ�H�!�@XTJ7�t�����F�S��y5����zS�*�X�rF;K��YֳGQ�B��/~ἳ�*�<����o�i�'ΐ9P����VF���$ސ�Qw��Lf�Ug&_	=V�)BO����#I&|��=<gRVAָDs���>q#|7�p�C�G���p���Kr`NMj�{n���p�
ݨ�<�\u��9�3�у�o����\�\S��:�]�stg�Y@�ÿ"���I?���k����T���$[���g��1��va�YKH���Y|��� ���3,�K�f�j���n�tGK�����(LK���=B��L�~2�+T��aO�����d��Ф�tiՍ���z
��L<?���~�LS�/��F::lC������gAc� ���)����^A�-�T>�T��&/=�E�,4�kySD�s��1����n�\xz�s]��Pؓ��\F�Q		D��r�ɐ4
N��]�["Bf����s1�T��ع;FSf������ۅɳ�B'�ߑ�c��l�9m�tY�{e}6o�e��$�J�_�+���B]h��*�"��E�C��/B9@мo���)�to�Pc�A-�����A�f�)Rhg���b�]�s���9.n���_'~��\t�(@�U�Mu��H	/o}�I���|E=��'��_xD%�t�3�WAsO�Z��z�3ƹ�v�in�=�ئtQ�@� ��g�Bi�rhYz��<�B���ғ���
$%�Op��L@��?w��Zc����:v��s���12�|�WO!��٘m�`F7�C��E�#�쬐V�ƔK��5��V���LlXW^���k�sWu�$	�}GCI�'��ejn�����i��M���)p��*�_Mz_�\��^u?�9����]�|{|"Ym"F�Y��+�h�=�Kz;�,n��\�䒲,¥�>[��>Cp�_Θ�#BH͡rM��)��D
2��s��I&�uD#$��M.�c"/�㽉���u_�̞�p� b�	�|��l��!�M�sNv��^,�1t:�{���yX��{dM��������J��7W�W�Q��G�$�O؁�5�p�Z�5W�EPgE���$Q�BM��]�~�#���6@A�D-����?��6�9��QFSIL@�L�k2����q���X��*��]h���zf��}!`�B�lA�l�\�adtf,��m
�@��u��]]�ヹ��#_��&"[���p�f������=�X�"�p..?g�yln�M�̐#Qa�
c��OJ�̀�<��ϻ�9	/E.�"I��#~�Si�\d��e
�]���I�X���f]�|(z�/G�y������nSG@�a���ۙ�P��@B�5����Lj���?l����t{�:vc�ջt��"�DI�n�����uL���)_� F����\)̣���ZB���Wea �$EG�7ܟ�H���y���{� +�~�!�5���g���@��guy�	�� DA܏%�M1l��ϫM�$��sI�>�綎\�˾��z$���1Z����)�Kk���2�`�q-݀�`.�@s�1<���3���'��2b���ݏJv�Pe{cОΒ���|�zR���2#���F5w�rE��-�D϶_�c�8@k��N��$Q�.EG���p�͓ygV�&_�`��%�Hְ�;��uAz�T�eΨp-P�`�HJ�*}
ۭ�>2�~)U�<!/�h�Qз]vJ����)�`���T�/�|9�����x�@�u/-@YC0)d a&���J��ɂ�a�~�9P�O�Z�}t��RI�"�YU�{3>"]�po��B�49��� VZ��OuiO*h?]p�C�jU�,����z96��>�|�}0�zY����ږ0Y�(���t�����4DA�1S�7����"[	< ֥�����B��48�\�^�,#w۸a�)rп�����P8�D7A)
�z�>�z���Sm-���D~��M�9����{$��x>z��x�ȖW����-ہtE_�qkef��O���S��
�?�oʻ,�Ȑ2n��إC��p���u؏<馏�z%Գw�L�ɱ\���ė�HN���k�����~�J�=�y?\�=5�f\��S�Ӂ:�/��D���5達]���?t"�J��ߒ�Y�J���r閖�~`����G>{��.!�Vә���P�L>{_/]ؓ��ǡˌ��gǥ�:�����0wQAU0'�N5���p@��o;I3\U��p  l�b\��0p�#��MP��^8=�&էp��\��X�һґ\W���$u�H���sH\<V���\g\���I�<Ct�I䔆����k0T��] uy�V�޴ذ� 5�/.EZ�lCm�A㼱1k��s)���O��vm�8«#3��y�M4�m�rH�h73������|��D4{<��?��XH���y�ƽ�Ο�Ѥ���@���=U������+�j�^���*�c��3_e�Ϸ鬌8!�zbz�O9
�=XZ��O�0�|#CƋ�	���)5� ��gd'}7w�M�W�v�r�'�I��Q'���5	ʳS�Fw	ȪV<':��Ǌ�\�]?1�ZG�LO���!�Af��̳=%�,6A�m�M�G�wk�� �K��l�;�P<�x�r{o/�jU�����+��ȷ���ʿb��'{ºmU�\�Hl̯i�N��k=l�,��ؠg3�����B��(u~|t��c!�E$t�3⒱e]<��� 9m��-=�

l��ڿ���m�C$#U�-��ȩK�ը���M����W�n9)�����<G�Z;n��a7O"#�\O�m&�DM]�=r�7�֦�} ��4��X����2߫8~����N�-���D��4{�n����R����d`���=:��s�n��ϡ��~���B%��i�t�T�l����xcC�Y6
Wl��G?@�yۭ	贐��D���r��E�����Ȳ���:��8�����P��o�ʾ�\f �>h)��[T���I��04DR�f6��{�S�W��%8����PԏG|�8J�G4�P,� �59��ؽj��cH�p�_h-�t�i���$����l�m$�����Z�^�Y��Ԧ-a��[�rexڧ�-� ����b%¿���	�:~]vA��笽�`�^�����nt���U���B	�����;\������d�%���;~�\|w
c�)อ#�K�>F��[q�Rz���^o�j~Jǻ�iA�B��,C�����,"�AM�F�v9���I� E�"�o�5{�s]���p���=A8 �#ɡn=�N尩��P�s&P��j6�I��dyG?A2��g�q�މ��0b��ނ���r���&#�i^��#99�8姶����� {5��G�TqdD��"vD��R6H�g�O:�l�_�]���`�u�X۶	?b�s�ϯ@����mI�|�7iO2؃�dC�V d��Ks��;�d�u��_%ʪI[n��I1�UC�m�7�t�"�%z��3&H�#��܌J����;�x�ϓԦ����c��ª0���邒S�qd�LO�&S�S���/����.�����39Q_a�|�UΘm2�ړC��/��7�	���!�F�$�d����씛H�T��2�=53�.���5�����ǧ}�3x h#�\��Q$?�=�Z���X	j9���t[-@4z�3X�{�OF�׶�>8H��}'��#~_����ޅxE�e@;����N�싴sjA��.���K۔�N�W��Jj6-8���#l���ӂ iј��i�������3�����ҧr,���(���w��v)g�Z���84�vJ΁�d0�3�Bb �����s��u���ۋ�Tr����w[�]"	�eDq},*�>��eft]��i�M�Tc��@����<�Z-f�����}n&�[��a��iRFTH�(���!b����PRF8Z�F�`��JuUs�KzB��3j������oPY�8�	��Dha��_2�ݴF7��'J���R{l<�DR��.��K}Rp��4R����*M����r�w�M�'�"�|ئQ�ަ}�#�^}��x�`8xN�$�Q$F���h�3�Y���>����O�ゖ��}z	jQ&�G�Y8�&X2]|J^9f^U^�w	
e�o}�5d}M�0��b.��u=�s��aԼ������Q�\���Aq��%�Y�O���<�L�G�?l�+�k&�2Ǯ|��B��;��о���{�)��Er^�Q����|7�"׀� ��y���2B$Bj���/Z{p4_y6�a�R�=p�z%�!�(c?�;�ޔ�hۖ�[Pl� D]�@s8�AƱ!�g�~N:e3���O$�)V��a*�;\D���C���LMS�o����/���oC��,�}
$��M�;y%|��5�z��AX�>�g���A�P�ri�?80g���Ǆz<�5�YY� ?�������t������>�]�Zs'�ڠy`�eɤ�J`S��Γc�I�őitU�S��>�'dxU���N�գ���ck�C/EԵ;�Gf
J���7�[_����\�!u6�Df���F�����	����	_��nF��	*� �|o�
�3Ey�F��h��E9Dr�	z&@�e¿��$
�L���c,�f��� HAr�1kz'�q�~k-��R�������U��n%�F�
(��؏��\��-6��{��:�KOBz�:QlE�I�/����WT��,گ�wW�/7�l����o):yo3Ǐ�Y����s��hT�1�����h�]��"/�m�?Q�L=z&�'ޘ����}t��=z�O����&����<5�[/�*F��w}8x��M�=�)<�`�s��ң޻R��z��o� (���.}:bQ E�J~��>%|�M�\�ʀ���G��/i��J��32��!�3/�\��$ ���nX�4r��/\���D%]��g]k���:�N��PF΀�U�7�{��Ky?t��>���E��Y�۝��J� -����k#.9癮��V>�ڒ����#�<�������൶�4������=�,4<�;���#wy.��e+�)���H�$�(1��:�mi����f*�H���軁O�
ֺ��!f�����dq;S��ݗEi	����?�e����0���B2T�9<�&U�%6��{I���4;�(�FZ�/��0��<,@K�KCRi@�<N�C����o���/���.�)R��\��q�JH��:I��4B�[ ��~j+;�c�qQw<uH�͋'xd��,]�M%�ԭ#��TN� ���~���`7ce�1W,pw�/1c�{�}��\{�3@d,��l��o*B1�R2��&��<@҇�m��RN��!{�i�y���x=����o�g���v�ۄ$@ݕ(� n�u��_堉ں�{�̓R<�r�<�z�C%���:u޸�6=
#��/\sI��'R_�����L��vL(�[[
Ds�@�*m!O6�HZ�^��ANe��Y.(=�M{���88�m8M���*0o��D���L^���a��QgR�]��#Ē#�Y��P�%M]�����Ů�II�N�$�`f�O1Yq��*=���frl���Na�S�zS�Y1���yHi2s;o�ګkv��W���z�1ӆ[w�=�q�𻺕IM�|�;Y�Ц�i��9��S��U0�>��a�dĘ�p0ߣn�v���)�jL�3�EW8�����V�l�신�5`���{�X�~Ux�N?�������Vd��W�����o�iv3��Ӂ��Ĝk'_!��u�@M��ԩ�����J�Y�H� ���9�UY*�tB���@	F�$ ai�]X��q���'���Ez��Lc�Y��>�:�_>ӆ ��I5,"gFQ� �v�zz8J�!����q�R�4龛-����rC�"���K���"�}��ܸ}{�~*���P��:�A)��w�9���TV�=�n�5�xz�������T�	�tm�w�|&�t܈�@��6P��f�b^�Q�<��Sk���ї�M���u��L���� ֿ�1Ky�� ���K�Ր}��q� ����!��O��j�l���bH�q��'(�X"�v�%[��?�R쯴BL[ qQڒ��ܚ����EP�����H�Q����d��ns�����
���	� ���D��*~��q�q~ـ?kZ��>YWم���#��Fd�*E:e�Pr���!G�ۚJe9VN���z�ԫm����LIQJ|�Y��h�
&G�'Af{�K)}��&ԗS�p#;YŔ�hXFǶt[�6��Z���C՟Vo	�U}�3�+v�EF��z� /��x��C����Ҝr�7��϶�Ϡ�T�9��2�@4~�����竣��P�Fz/�$����9(V�
ߏ����X=��}>b���tH��=ַ�#E�
�C�CLͼzy�5�ZH�f�n���܌3���	�Np'Eu���L��iE0�,�º�Ѓ�7Ȯ�}KH����`���M�r1.�/D�$i��W�`렖6����*;�^��ԟ���U������be_�(�u������Ԗ�+�����l�]>��dZ/r� �0�y��=��d���Y麒��&;���Je$Q�甊��B���T���������jp"��':���6������`��������N	��'o���$n7	�d9�d�`
/�ϣ�K�hK���`p��,�@W�o�D-(�5�C��ck��ֲ}�����>���<�gċ���F<"a=�c��&���o}���E�r�r��X�������g��
�=1��&Aޕq�Z�nο�<S�@M���H#���2%��@`��Q���1fd+�0zb�L���~1�����u+t^ ���L�K6�*�m�_{ź�+�﵋̣���G>���D���
0�y��}�ō����a�N�a��o�7��!��Ifʆ`y=��}�Yl��p��r���Cd[���G���1+D�s�� aAa���ؿ�x8�+Zuղ_n�P�����i7]�L,gB��N{��-�[�0���D��[K�ԭT�O�#��(�-���([n��Mr�5W�K|z�j����謮Wր�qa�g�5�(��S2�`@�����hR������4)��:x���l{J��W���~i+�lIf�\c��LC�9n��x���+�����a�|�A���o���?�ȃ���jѼc�Zb������0�R7*�<g�!��dTyY���Ƞ�i�wje���ob��}����K8t����/��ѯ�+��[���)"�r����k���Ι[���O�P�V�1�_���w���1� �R:i��Ʒ=N��8�I����J��*J��E�8���`~�d� �;��v�ѯ��v9u-��2�2v+�S��y`MC4���@��*�k�Z]|����O�N���$ƭ(#��O�ML�����!��n���;L�� (z� v��1kL��q$�R����,�$Mb����,����i/�3e�!��b�!K&�OM_0�*�BoF�29��n!A��z�z�D|���-�DI������.?u���������D�i������{����-5N3;s�����o	9�ժ��g��h\����jv�&�Q��R�E� Io�R:Ww�p4��J��E��G���-l�'����Z"� �0�{������fl�B��}"l��X��97�# �my A��a1m(��SG<����J�}��wFo��T1��{'�۷�	��SB��W�I�W��=��(m=�� ���^5*b�a�m��g:$<Ӊ�h��k�����������5*{a_�(C'G��f����NLXo���E,Bl;���a�&�D���TA�i*��,>��ߟ�$�	r�c��	�3�xR�����-QSkf��K
H�A���Q�
��ci�K(�+.�[���4�{��hCeP�>ӫ��O�o?Xu1^�_��|y�<3-x��a�dTbk��i�������+HF����ۑ�ĥ�S�~�X+�����r�A�ƃ�Ia΁ُ�e�B��=�uk�[G.��F�W6�3�0L"b׊h�q�䑉u���+opp��1���
�H��R40[��Gh��쟋�%O���_Fab����:<b��q*��R���U�g��q�c���uŮ�ad��:�k�F�������v�G#r >D9�P�a��$�c����u��7ߎG=��E+�ӄ�Gc�{���A62�ێ�*�VY�����d�_����\�p$j�P?�K��G��Χ/��YX�S�����ޓ��z��h��5jYS����Y5l$�2]ēJq1L �r�ӄ�p 0JK�Z܆fD�y/,��r�T�_�R��8����&T�`o�Pq��u%�/� Bs�M�a|�<�Ha��h�ZU���&��h��M�����Z5�HQѷ�4�{�-A6�]瀰�B�LZ�\ p����r9��Kj@�J�9��5%�������!�0�㋿�9��) ��J�k�'5dD�L�m�eu��0X�6Qo}�D�˩T�Qe� @I�7fF�R����rW�� ���w*%&bݚՄQ~��Q�2�����&�%��9��~�VB������a`�FD�����}�0���A2 �]dn����J��<tP>�*����	���>����h�kz����9�*��ߔ'r��蝳\��`��{��Ɣ����ϭ���v� ��L��X�����6y�u��M�����G��9������®� ������9��6��Z�e�(�G��:)��R[��ϛ.�*
)����-����#��>�0d����o���S��c˞a�B���P�s��#���f�6���^��|6�RUǂ7�@kM�/�=+����(�1%'�e�`�-R�/#��ʾ�4S�R0�g�L\uɣY�x�ei�WV'}uŎA:�_�u�8/DWJ�=�e���jR�x�X��i��OB+�DV����Je���TC�������m�o�;��̩u?��d�c`΀��_�㽦z�k�qM�P�(Ք2��H-���`��٤	�1�;ݏD�>���>"fp�����^	�:?`#q~�h�#l.��=�S��BIP_,0�
:��R�g*�S���G�@�֐�mΕJ�c��yX�s��X�Lc5��b}'��to;z3�on�� ���7����)�s
�P��R���gl������#��+��l��r�8Q��ٵ%6Gܼ?�K,/-��c�����Ѕ	�v��AB�c���9F�G�u���)����>��ii8׬#��`8�%C� ��,�_��
��f*`*���������A-�5<}0��(�^���$�/�)F�>�K��zkss���*D}��k�1A��~�,Q6��>�0�}�-qǅ��V�Dk���`M�I�O�J�2�w�I(h��K_eg��Q5uɲb;qɵ��IפB.�G4�o*�:bEL�[��2�O=�66�SA�z;+����O�}T��X�ܓ{�ë�-��U��,�����s��1�l߼4�h[N��M��a�C�D�Y�]��.��&���
���y8o�;wT8)��W0��ҽZ�W��͊�k��v�g�o����F����'^AikE�;'�&�AE�hLJ�i�1�I��:ն��h${\��<�-a��JJMG���A������S�� ��]�|�\_ϋ9�8o[�i�h,�n���gT�B�T��6( *]�rz�R�navSR�ې��$�o)�C���Xe�&�x�ev��N��q��@<,#T�$�;�+sO,<<�/�A��ڲ�"J��T��K�EFZ�t���`������N�Qܲ[*����H�w�3����e˙�s�_KKT��^ �t�Sk�^�0:aE��F��l"��+�?|i�y+�̩:�WSy��&��\u������|�>�f`@������A̠�3Ur'\�N�����뵱�<wa"�Qg�JB�(@�Y����P��zeq�М�Z������#ڤz�P��p�4S�(h���u�4��uz*ׯ:\�ebp���?e(�yͣ8�U�b�g���dj7 �˪mʶ�I?|sd����%6Gk��	
G�U����.�6N������� ��?b�ML2��Ro�=��+�C�-��5=`{e��R��F0���`b��됹r��v�9�9?&�U�,i������a��r���o͖<����[�@�z�/�|�a =�8�࿫������г����Ι�ˡ_5�<t[VIf��w��X�
�ujE!������ؕZ>%.�o�⧄��SY,�P%D�����rՙ�4��э}��Gr��ka�K'e�ڸ��C�)� c)�\=�f�������nߜ�-�u�iv,.k���l��3�/T��3�j�oi$��1�ü��j�G�qli�I��+�b�x�]�����p��v�z��&·����j�llVK��IS�~b���k��N��~���q>�ԩ&��#UW��?���@1�M�37�u ��`dSz=��+؇��=���X.�b7�$�c�;��Nnm��	�b�\� $I\X�l\'���O�ҬP|���!(?�I_�}�g�)�ի����B;��wN5�־S`7Q⒗��JY#���au�,��k��9��B�9�FSձ�8	֖�Ѫ�n�a�VC��y��ćV��;	��1e�e�ѭݳ���T\/5�N��&ё�\_)o�b4��ۼ�t����S�&*"F�e�b�&Ӡ4���>���mm>��4�c>������ꦪ���t�Ü����3���V��F:�{�۲�m��l���m?��U�J�K��U��B�o�1K���븞&k��x;�H#��$Qh^_��U�ef��٬{a��^Y�E ܌=-�"�Rq�RM�*�}���2��L�����z�?P��88�2�A�����ۣ���֑gA��&4�9�E20
�y1��k�STm&��dwK��H\_4�]$o���VP챶�Ky�&f��V���q	���`&���tM¹��������J���+�2�ҷ�z���qKjC���)4�P��ưv�Yp�c+�f�&�ѕ��, �Ҿ�A���.-B��!}œ-	�a��d۟|���]GN'5ƭ)
�7$�J)��N9�͒�I�f2 zg�۱�q\9Y�{/�H1~�^�x4H���%�.�)����9y>�T`w��3�f]m�h�^��o��j����I�Y�U�:&H�$�#3�����UcT�ƾ-"J�I |MJ��.����Cѳ=	Zf��8v�k��u�̡�ȫP��2��U~-�.^�"W�D� �S |�A,c�lx�������~�#�G�8OaP����h�470GPr%fS?�y1�VDN�!(���z��J��e�$�H4�%owê�kjr9�5%��w���-�J��A�9���a����C��.�1��$���*k7���a���8:>޽�����h�|j|��8C�0������W���ːq *�=�����+f�)��#��53��D��2�"� 3�gH�9'2���sJh�Y�"�_�f�����Qi3�w~�����ZG�3��}|�T�� $��B#���*=�6��&��`��n������c�;̴��p���?]pj�i�pg"R� ��?7��®u�GB��DO�ߤ����z;���m��_���++c��=�TB��W�'�9�y�����' ZUV���0;�XtST����|�[Jt�S�dZҾ�; ��`jSlM���qJ������Z�Sf�x�y��Ǒ�v$�EE��&p�Ҩ;�����1���|�&�Z�;X�����K���ZT�����%,H�v@���o_��ज़P�5��l�׫���΍���z�[vFXܜ����U�����:��ވ߬|F(���P��j��:�r���}H�Q3aQ�d���ݢ��T��Q�1��R�8#�n�a4��)�++'E*x����V�F0��	/����^�!���s��tI��^v*�!4���gJ��3�?)ҵ�pf�%Db{��a@�M����e�~zZO���/ ��*>��?���2Z�C�_M�3t	��[2k�=���cm�d���K/D?�8S���)aA~�T/��	��J3��jf�9�}���I� ]O�*6g�5-��nݗ��9�ޝ3qˏEX��`@�Ԫ��v2��^�;p�K���u�� �Qo���L��:�L�u|��;�GX*���~Ne�� ۠���s��(��b*$3��u7r�t��p��,�%���:�����uS~7Fnl�Ob`���'� Z�<:��Uz���xu�%d�4�Ȃ� �Z1����UfעA�w<?�<�P�ePT E���N4J*� "�[5�/����1�5h��
�C��Sb�6��\\e�.����Bi�+5~hPai�&�n��Wm���'!m��Ө�RV��\>/J�ll,OS��<��ڌ_5RQ���Z$-Em�A(qo��sYL^�&��Q`�k�u+�M-�^	N���g�^��W�Q1��UE4X����K`�P�^!��Q�6>c�5~�TF�c��ٟ���jN�;c�yG3�gZ|Q�R��l������!���sS��Xg���;p!�@���l_�6��W��E��pDQ:sB�JCq��3I>��)דOY�`�rM� 	����s��tq��� WjO��J��z-���i��q��{Q����G�.�
���+<�B�����]������i{&����]c��V���E�����X�g�c�PĚ��1/*�Y�����p���4���ޘն��MS{���^[�3eY��d�hS���2t�?>�y�>�n�J�qN���AsG�s��UW)�t�U��U��m�g���!3�x��żܓ�bee��
��M�T��ȡ^d�_T>6%�1�9h?nu�Pi,$��L�J#K��j�1Ʃ��^���[X���ܝ�� �L;&�V}��O���K��؉��(b�[F��E�q�lH���c�;]B�mY�� I�7���1ZZp��������v��>��S��6*ϮX�i�r͔�(�F\?oԎ���g����~�Pȃ�9+�,`��qU�awS0Jny��[RT�N�֨����Iw6�����-�����FVt�R�|%W+�W�"�U2lq���U�u��&|J��7X2bb��聱B$V�me��Z���:���qK�(�!!��E�؈.Iޚ��ȺL�	�
pqk���	WL9�n�}�^���64ȿ/������6s;�>ƪӨb 1x�M�f7����� ����Jxe1�Ͽ�
L�'�͍�є�B�X�SƇzK��C���/Y��a���o�J=+��qh�/��Z�'l��nlm���3(iӴ�ǥ=��<{���Zߨ��U��Ϻ\O��`G�;On*
��'�4�u��.X��C>_ٗORb%����8@������:�C��;F�#/�V��b� ��o��l�t�����;��R�0*�P��2&�����N���hk<�>d�������� ���1��Gk�iHY�{B�9�����6���3,��F�c6����IvY�t���%�䛎��Sk(�L�sv���L���dR�C%�ưY�7�Q�4�l��Wy�k�� gT ����v��|����I6[8�t�pt���ޢ�'	�z�֦B�Q���O��E�K�h�;' )Ð'o�n~:�Qj7�"I��>��j|�Gg~��s	7Pi��J�}7��e���xK��w�R�}V��آ�>(/���\�rg�>���v��f�ݧ�{�m�L+������If���ZSԄ�4饢py0	��
�72]Y���8Y,%p�hwg"�}���h����|M*Q����=5[jTI�H��`zZU^(8�x
q��rRg��D��J��q� ��l��J�Uu�y��wH�ء��h���Y0F��T���#7!B�@��{k���$�g[>‿�@��<K'z�S��0jL�;`=k�H#��~Jl�ͦXp�ч�\�į���#��/2�*�n�Wm�򇅸]�k`QZ�{NL$T��D�Of�&��:H�*�C�!�Is��I�W{Z�J*��-|4ϳ)�fxY��f���{���X����Z�_�
F��d�~z���N�;����Uz�9F����U_qU�:�ӓuL��ڑFL %o�~���0�\t�{���|悰h
�m	�m_U�2w���8��$���L�i_F����`0~��#�#�+$�2�K��#��$���a��{�k����w�a�z=)�g:;E�	w��~]�`N�SU�L�>Bwb)wa�d;��wv�x�T�X$�Ȱ%Q�b���5�J�i�r��b�/L���4T�L�J?��9է�ݙ3V#R��4CMI�?� Mt�ZU�pL
��s�c���`]��ɓ} %�򱢪���G��\@���d���s_E@�hB~ �k�rB"�)?���`|�15֭zS����� �9�nm
&<4�_�L"�Qre�q��	F��׋Ⱥ���YG4o��V��f�1ԗ���(^�Jh�Ҭ-#��v��mX"����.�AUss*b>�s�@V�)x��tI۔�������'#�XC�o��� c�؇�	,H]��[�$���ڇً`�1�j�ṷ*89օ�����i�}��T
G�j�����3�=���m�W�w��K�{bu���;a��N����e�B��e��i�í��Ō7}C�v>{�&`޲��n��.r[-'?8"-n�2��!K��k���|�+z�fM�`�Z]d	R�a3V;H6a��V��R��xoC�	Y:l����XyGI�T�y�k���+s�\wz�oK �jI����>���=d�sů�=�Xv�=�`"q�O�A��o�-��)�N��4_����y�$���+��/t8Wu�t;�j�e��W��=�<��2x����<@ -�������d�h�_����~�q��N�C{d$�SBB�����[�E|f��ƦW[\�����ri����>��,3<�c/�T&���I�Q�I�S[s%�h�|&K���+��S�Zy�۾�-�4�Țr߿���lGv&"q���b�1'=�w#�O�y��t=��m�l�IqUv��I��J$(t5���X��%
m�ܿ�O�O����~�$�S��F�^_ǒ�A���j���.w�|������#�9��j7H���)�����
j���EG� (	3�'�tf;�Xh���]�h�la���0������y�-���'I:D���a.�}�0�z�����8�'������tz؛���cC���Z�i��K<zEG��beEX���?Z�u�g�c���c����7t����wH�.6@���O���kKf�f����4
�x��R;�}�r�*@��6)Wz�)H��{�R41%�\4��gR��'/T�@NC�f��:̻�iy���Q�9������b�E"?��|2��zY�ք�1�}����]��	>�~�ɧ�S<h>l�V �����3lo6��OUL�E�2�U~�� x��t���XroD�(`��~:�O��A�ܵXk�u0ɽ�ЊP ��� t�.�Ky��v�#���3��\��)	�-ф�� ���O\
ۣ�y7�l�C^����!�6�Ϯ�#�_�쎖@!]T�%9�����'�SW?sөUm�ܘ��<g:��{�+Y9n������Q��pLc?��ـ�Rzq�Zj]#�#���h��ؕ�jWY1;��A���^R�C����SX���{���N�뒔��p��r�`UՓ��']��cܜE���!:�ܹm%��Ɖ�`'��.?s��T=c��-.�r� ����&��+�O;R�/!�4Y����H9��Sv�"��s�^��/X�SB�*�-֮�P��"H� L���G��S�3�{�b�8��:m�8p��s�����Q�mUE����X��{6Sn� ���e����٢�	K4�g��$�k5��d�H����G��O��Ume�n�,YV���q.�-���o����]4��0i���T%��f~��:�2Д���Z@�1��
�ͻ�[�����E�H2���?�2�>��{��ts�Ȍ�k�L�����Dp��9��v���*������ �w�=����s�u�`�c��n�-�-i�:S��d��>���ݧ��rLT���u�z�Hyp��	��q��,���̜���!g�"�:�c���˰�H
����gG�j��50Y�K�������OCɱ���۲R�T�Q�HB��>8��O~�#5�!�ZBG%j�`=`)E����3��R��1��� �&j ������%���uJ?sQ��4�����l�����/��U1�_RW�?��?i�}��d�:��)_���.R�.�+׽�%ɆA�`o��}4@?Ŏ�)�5ͱ��xV�{���Eq��C>����@ø@O'�����Rz�ިU��U>�Dc���9q_�{xD���@��Ö ��waٸF<�T�U��@�m�r՝�[Ӈc������mA`������!�MG��P��W��u��}	9ЈÌ���{�#Y�G��%Ӷ�@����aEE��}3e�U��@O��R��o�-K��������r�+`�섲��C��2M!D��j�~�0�y��o.������@�Ѐ������	�W����=����\/*����+�˳�GK�/2ά넉���H�?����'SH�wBڛ�sc;�)#���aRhV�t��������Iž`���Z��
��oƜ��]W��x}z�a�A���q�D%B�1g������WSZg�S�R�QWL���5#_D�h���Y��eŷ�:�}	;��.A<���ȭ�t��H�V���>������A��/��v������]S7c��ϙ�,4��$�t=�6���kE��E��v�B���M�ӮKs��$ G���'�ݺ�,�cck�_�۩�E�n6ǡD�݋+�v�-bqX�%�I@V]����I\�.N���_�TUH@�N��?*�u ��K�˚:���%��N��N:�6�y��t��@q�q��ǈ�+�3�&�7�ܳ��-��:!v���	�V3�yɒ*��i>q��I\�����/Sy���6��-���|ݾ���$C#�E\�t��KO�p�$��@b�m�[_�O-��?08��U"5%��)=��`��Ʉ�k�Lz��I�,�#" ���h�]���Ki��ask-��:|����r� �7Q��
#�]�ܘ���I��f�4�Ϲ�����6� G;��"r����2׳�? �1����N�i\6�?���ܦkAL_ךQQ���KVh���3��[��Eн˼q�@�U�3�>0�0-P
��,GMYk��V�dΝ����4x�=��A�P#��;��S�y��K�!W^��|a[�?�>�;�Ĕ��v�U��~ڵ�˩��.h�FLw��y�
j>�\��ID���ܬd>�-~�gf��H�$8���4�.��a)�U�����
�r�M,���kA�(I�q}�O�.8bEʅ7e@ X�۷'�'cG�]@<��ߤ�n����"�#�;�y�{)yK*;�zGuO�w��K�3�p���_e٩S������8[!��Ge�"�f5PL���TO\z�����63�nh-�^ rO'��M$`R�)M��a��܎`ºNL���PCBx���
��!�K��N�!��g�֣w������c��kl[FY�	��}J�q�3�-O�ѥ슣�t}�.:w�k�4���v�+H0�������k\�"����嗇à9L�4D(�JАX��WLy���y�Čs�t����^	�U�=y��b����v0����@^"�<h��7Н��':ӫ5�+�1�dv	hi�
��̉{3���r��X�ê���b %�w���E�đy����Al�c��!0�ois�M����U�p��t��iM��Rvo����p�L&S��͖<���:�Yr�A��ϫ�Q@�?����h�I�P��0G�y��d+l$��$���ͅ�T�&�u��h.�K\�[UbQ��f-�:q�+1��h�3�'i� ���_�y��b��k���4�����b���Od}�u�Z�0I���b4�Q���O!#7+z�ȓ3N#{	q1��T�ВW�G�ΐ²g5����׍��ܗ]d,H_��:lP�v��H.C<ϵ��d(��2�(�-{o�����������ˍ��2X�J�5�߰��Gb�Ș@��4��C��g]����4��[S�C�����ɸ~��qN�(���y.72�V���pI�L �/�yN�U9��9��
\j���U����l#�5*���[IK:Z��{�3k�ۃFk\�d��t���k�|��(g�3B����G�~;�ҋ;�����=�񭦧�1,~O�@+�N��u�r�^O��u'K��R ��;�z��0��ǯ� ��*2�2�	qV$'$�/�(�0���#U�M��K�}�����d_�T*��sr�$0��bDDα6M~ܮ��9b������Q��riA���q5¬F�m�s��Z�֖a��sy %ln��-~�*����E����S�Yv�g�i��:�x�ߔ&�_T�����T��h;5G7��b��U�'�@j��}Q��F<�&���� ���Q�W�<3���(z�EY����G��.	<
1�c�_�l��CW�� �Ry~�7���te�2�C�B;�B�Oϵ$��3������eXY"҉��m,�7m%�g_0�K;8��r�>�d+��������H��x@`L&�_3�|Z2S[1#�9�6U�k�"�c�nO�3�͕w*<o&3ZI���u�����BG�]���߽qM�"茽�1d�v�<�m�oMw�0���Z��.h�2�j�����_��'1ķ�@j~�h���*��8��;����}�j�
�Ϙ�y�_�n����Y�(̄1?���G���Ox��O�W���^�b*,r�8{��y�����L�h�P�5�bv� +e<�-�"w���Ï��F	Og�P�řz�Xp�/�fr�7iA�UDm��x ^�/]����A�fB4�Nht��l�����7�(���mY|a�������_����7v�?�p�������
&�=��Sz��FB����U]i�ȑO5��Y�?������<g)��XT�&�N�GE���A�zE���*�e=���\r2�7��%'���|��)p"�W�,;��SĄc��0���f��ف�-���x�KfI�\�8��T�y�uXj8h(���#��G�^�4>���-��/S5�b4θ�h<`u�Oڃ�Ǳ��)1s��o�_1NrIo)8����:`!�W��7��<pCA�BG>vD�<��r��$��Х^{��G����8��AV��Eґ�:h�bOe�g$�v�}8m
߂ý���@a������k=`&vV�'(ӈ%�]ν{ʽf7�s�$�����5(g�]$U{��-Jw�n ���j�ɂQ_m�2���+L��,���(�)�3��|�n����?��x��u�B�iA6gS"����q��b��H�v�A���<�	���]1�b-Q�+�#qV�b�BM��#�?؜y�M�<�����A<��|���n��1'��88�˚J����?TA��]k�.[I�"x%&"��	���{N��Ϊf���t�W�1,("�;0�����u�Cr�uӞ=�s����v�NH�.R�!�(���̬�Gz<-W��mI�ح��=������B�da�F��C�`>/o�� �ˌ�P�`�j>��E8l3��4�v�����P�z��#+���([Њ�|�w�� �f_�}��5(�[<�]6Cꤗ��GB�m\��я��=�M���,
�}Ev�ع$M��� o�un�c���\I^k���\�xF`	1�cl�7~��>K�~:(�P�ir�Ʀ�����@����֚���??tckX���g��y�sx چ���2=��C�����]I��A%#�+��M��ht2�%�ǿ8��!X�����z�ľ���^��C����A��P��
�ގ�.5�� }Q�����.A�p���4E�@�u�^ �%خC� p�_��Fx͕��#P@�_����Ӎ�ӿ� �H���P��=��J�����G{�	�����FK�.OU���y܎Ta!�5+nP��Ts�TFnCU��,K�U���A𝤒(r��:�N�X����t�'�Y�Q�
o}�����, ?�Χ�ƕ��	e�;7c�l׆��r�%��6/+�����f�{��e\u�+�>�\��z3�
WjW׍�w�p�u��G�����:ŭ!
CJm�e2py��=��&}��,����u7�X��I�9Cwpq����[i��5�.��]=����.�i���ϜB�cm�k*-X�^�}e�c���ƌb�&o0y����WW�=�96M>�
:[�p��̬��Mw���3�Ks��8	�¨�A�H�ԐS����j�?eH�`���ͼ�FN���T�7
���� �1�)��^��Τ��m�y]���S0����=��H�D�W��)-�Z9�)U�$��^�������n�!u��"�?ߺ8��\@�5�'�)���i^�n�$��!�s��VuB����ĳ��	Ƨ��-��;:.�KZw���L:/��X����z��e�*ȋV-C(5�oB��6��/�|!���=J�� ��6`��G���g��κH����K�e��qJ�D��u��Mr��UR��E�Y��Z%�G���"ϙ�ILk)��lϤ�np��X��[��x���$��ڭ�a�]�v��f��o_��L���GC���L�^%�ApN�G�nm����f4�K��Q[W��6Y/��ƊZF���V�
:��� ��09O�(������|��,��>[v{e# ƾAqjO-�+��&�?�2
���PY�N�nV<]��aĢG~�{�\��aP�6E<�_�J�}��a|��1�s�#ݽsG���nF��0�ek��~1�!c"<�8�����f�������B�J�'ʘ�9��G7���>��"�^� �"K=�XS�Ҧ�q]?T��t�r�V��/@��b#�\Ϧ�8u�	`}d��w�Q�)M5S�(2H��|�*n0O¹09,��l��،;Cp~>����(~���J������2>xE� V-����Z��,���e���`1��m��f�ۇ���A�VHa�_Sج��:�`s��2�*��c��=���������]�Я���s-5�6���e��ĿC9'\_2�Of:���MN�`3��'v3����5<��]$�)r�����o Q�sv��N���;�V<x�6��FMX�)qHE]"��
]�EpӞw�[���C��{��B,�f��։�*�s��
@>�?��ŵ&��2�kʩ�۶}T�E�zD�?����
{ǆ�s|�?���WnB�_8Z1�ɷ*�%��NL�uɭ)SƑM��wD�*��b�֭қ�
b����3��Zv�߅��k ���A��bP�D���<e����
$ֹ�|�g����Ϩ5i�A�!�_`�9�?f������lX'Ģ�@���6wv���f7� ?�T�Ƽ��)'"r}�o6�`Kg��ݙ�B`Ie� �}n�k~t����(��+?�e���Ȋ�9�������:o�K"ݭNwZ����@� ։�W�nc@4�2�0��,\{|�G��=�C���R�A�N�~��[`���J�)_RT����ۈu<� g���0'���ir0��]��^�R�1q�1�'OsKk�6��f�bې@'��\�d�p6;���q�p����V���<�sj��_���j�����jmz��<���� ;'�h�*���D�$&�a������Y�8�ݕ�4G���������c� �1z"\0S��Ĩ�DE��ͫ��/X���1YC�w�������2��)������l���v�D��N���R��w�m��Xbo�\rG��4��eo�>�{���:����Ɇ�M~�	�~�C韢\uNИI��i���חF��
^�V�[j�ob��ԉa����E�d��B��q���#0�%�'����)W_K�"�?4��'�^疎�@1�<�s��d&��b�g[����׌���P�>��/�����'Sڲ�����w��$V�>��������&�S.C5�Z[�p8�
'�8ܭ.�6 �()٨"烰�E�t�N���5�i�o�=ϓgB`Mg=��h�G���ʋ7�<��`/��1��6NC٢��ȱo�=�n�
�� .�h"�9���k"hk���,��(�W�{���Ԭ�7b#�����;P�_�w<ꄡ�Ϗ����s�����O(�����q�����e��X�t85�BEk聛�,\d�&e�m0שȈb������>��}�X7�f����Lj&S�#�/a�p��� $-�����N����d���+H�C�g7K�-8�Q�' ��/2i�%U���q�,����Icna8P#��"����Ye����%�cz��D�p2@ܼ��?�9�����}6�V#��2��jl��A`<�F��#���M�u��� v�~�� HYo~�0��y6���3u�f�UWDV<;qwd5K�@N(jY�4'5���V`����"�\r�Xi�CU`�}H9��� �X� �i,��`�e*��OQR=6�7�uVB����"�$���Ӈ���Y�3�(��`��P,��}Jv	0o����2�q��W��.>�e�ca�y�@�����Mt��ԧ��'%}�8阄5E!���t>����n�3���7O(�X�/���mh�dN�"�	���l8T�)U2Q�P����9��U�KQV��$�q��l�;Դ�Y��:+�ZG>j��ƕJ�+���ҝ�g�1 �
b}Yp�"��ʐK�«�j�L�٫j�P�#D��ft S=T��L���+���!g�`�T~��M'�h� Q��f�����J@H#G�qp_, a�|�̀n�(�+����c(�s���Wن	C�!<L��(�n����� l��ًY��|~%�����8Sl9�K�U���)l�|Rb>`�ͦ�m'hW?nҭ�2��ߴ�V�����������0�^a-�ݼ`����%�RLKJ�$(Ѹ zo�~$���z�ߖg���ZG�lx�6rQQ�ztNZ��F����7�Q� �o��@�ʻBMS�`B�~���)�k�ѲU]=T;$)x;Ul�`�d�k
�5�XvYV�C��@�[�>�w_t	f!��M���Gl��9� %��t\P��nU����cG���%�_mdD b0شc��Ap�y��+�꛱�.x�+�3%��i��ϕP�B�5����&ԆL��w�� �#��W�k/�(�.�	�n)��[HS�f��T�`m'abO� �WF�v�Dե�Q��ٻ��'&i���)���'�������b�r+�A䲦�@�F��J8�X�����h��2B��6��:��X��������k�!;�g���^�v�YP�f�`ކ���=Р+ߥ�HQM����}�E'�H8ɀH�J$���B���K�>CU�,�D�*Ѩ7��=�#{���@�l���/�o�S���Ŋ1��&�����_�s��o%��4(��I�����N�Pu��-�۞/�g-�m����@�˽�_#UX@��~�Q��G�k��N�6�o�x�	��x^���͊�"�85�^S;��/�Z�0Ȣ��Mܙ#��~�o+�^{�<�Zu����$�I$)�;D5Z_J���ԟ�_|�i)�%_oÕ��ڽ�շ��1қ�bnYQw�a�?[N+����'�K���m�l���<u�}��&���ؤ��U����Q��3<�(�M��B�wt�2?Y3P��䅩��Jv����r�YN�#+�L���Fˏ�I�?�ײj��n�]�,6S�\����Ͻ�?XNW9�4?�05���0��rery�>��SQ�7���K���?Mo�8����RZ���ǝ��O��r�y�Ŧ�N����:�WE3q�Z�q���Y����fi��(�eB>I&5����M$�k �}."wQN�̛���|x���n�[�K�W���n����z��?|3�osh��6��D���	Jc*I��s�vC�4�s�T6t�VK
��Wp/������X��E��6���_ �;@�¶?�cn����Yg����㭠�q fˋ&|'�Dk!hWhό�G��9eY�Yl�lH��nt5֭.K6q�&��d�DVRỿ�I�D�~.~�-s���T��##-)@[�g�QeE�;��R7�c�J��6y5�qq�_H^1�?�2��L����#S��7)�z���s�Z��p�w��M!�-��0�3�9��!�������������.���h� %�ȉ:sz�dr���9	ji��E5pgLK�.�RHs���i
1=���1��h�6��8G�N�6F��őz�$v�:E�@��9Ț0:%�ɶ�l��ᮗn�/�����3�����|j@���D���;�^7�5N^����m�o�9�5^u�}�a
��,}�: 9��8pj�Ґ)�<l��o`�"������Qӣ�X���f5>Ul��B;��^�_�l=j+�c��WY~j��^�(�N�������Fnd�+�a$!����\7�[v;�Z(_�c1ܟ��緭�T�K�9��ߝйX���g�C0�<��`���7�-��o�Ж��%hĲ��{nH�S�칶�5����ʒ>gU�g���]ؗ5�p/��iRi����ŬTR4E{hS���)�z8@�O~{����{�ۺs���t�p�B=��{��@�T��h���$��ա
��=O�bt�J�#`�S��a�憣��0��t�%�D�6=��ئT��9��>9�e� �3��ՑZg
����_OG�^�P�I>��%Q �cS�#gASpq�b��D��:KA�����li�9���뭃_w�a�~�^�����(͞x�?���M��E71�dew��i�ej~v���?��#���uM������Fd���O?��@�r� h���<�xN/�#��M�E�2���7�C0��o��<_e��O�iZ�5��ʟ� ���V]��+&cc�â�����U\>����s�����������8���c[��:=�EK�(���/-�� [z52Ǫ}���Ӵ��Rԓ���Iy��O-J<8^݃�rc�WH�Oň�_8�~9
�E6*�+�W-����np�5ڕ=u��%�u&p�iE>�NQ�a�)G�o�۰#��_1Oq��f��*�c������t7V(��I�fh�@��$z��>�炔~�@�̏>�^�;y%D���NCĹ�u�D쇳l�O�]��a�dV"�¤�8�gM�fz�����_Ƿ�xK���.〹ǰ��D��������c�>ߤ�a����0���D ȍ��_�x#���uX �j0�c���BrŒa[\��p*ɋw���no�r��� ��g*�i���V�|&ڇJ�Xw���e3�S��*������u�A�v�uR���৺vAH~���	 ܾ��EWtJ.��<6�R2=��XJA*U)ע��ѯ˂����q�G�����tɩ��COJ\bIo�{������?8>ٍ1B3#��%iO)�(ZU��A�u",~�pz]2���[�u,k[f�<���&��R=Z�_G(8p�4x��g��7�ʉwv��s;�}Q �Y�,�.�����1�9w��X�z�ݏx�����v��U�[+�^�x�[$��!䕠Ì������Ye�PQ,e���Ԇ,+)*�L����_���]wQ�E����%�UvY1����0F���d���"�H���Y~�W	�w���Bʳ,IY�E����4z��q\�|�|=i~�Na@�ȝHM`_D�qs��3ݎ�y�!���F��!����	���Eq�s������V����!����?���TV���YL0ܫ� �]p�zdj���;?ƈ���3��%�ϩ������DQ�N"�.�\�'���ul�-�D�C-����Z�U�\rGBi;hM�D3�u���-Rb��Gc�Jm����`�.Z�Aˣ-���)J�i&Ml�]����$���FlF��Z����\2'b�lċ���7*�H/�q!8���f�$~�oHuR5Y�>Zd����0����/ �E<���h��dw�puf�<xN2��.M���s����O>r�d��
�;�k���2�tUۜ��V�������`8A�Ivp�Ey�ہp�)� �:e2�Nf�^���-��CM�nu��Ftؚ��%�PY��8+��U���@�Ã1���/��0/"�z
f���������I���4�pA�"p�\���rE���^����b3r�_M/�n[*U��2� .%M��:3���l=Q6�x�F��.R?%�l �����Q�?�WC|I�d���fXzg�o�����H�Õ�����BO�������Uf3yW��_T��fTU�����	DW�SNU�4#H�JC ^Ō����91��F@�L�].QSA9����j�J�j4��e��g�C0�*|�ygر��).�\b�'��Qp�	ĳ��l�[J���o���Vm,t2��{ �^-��t`Gz�d�����f�8�װH��M�w� �d��qt���҆�O�ͺ27ߗv�21ZBG���ZT����z!������p^���X|zp5�S?Bn�_���:���糎|��i���T�e��O}ۃJ��|��,��%�@�z��,0��C`Z�V6��'��.�J:�Vo�s�?��7�\�jO1�y[��K�Vf��*~J�Ǟ��^mI��HksTeD�2�:x��z�.J�l��R��f?��o�p~?��rȴv<��e���઴Ř�-��Q�ǈq��W����J�Q��� ��P-�0>�`,���� �:@>��+:_�>��~9���{㎂�͚����K6 j�1�^V�:����\�/�Mu���[�rv����Z��o��S��aE����b��^9�}�1�u�T}��b�W.����1=G���苶 1��T/��C�Ȩ�CP	����;�2��;�9�`�5ۄ^/�_j�}c�K��z	����Nܰ���kv%�2���|�rT7{ߛ�+>ζ�><���	�w�j���U�!>�#��6x�9��� �9��ƧD���B?\n��5��Þx�t���c�X[�e0 ��h�CAu�6�j�mR%�B$��k,�����ܱ��V}Y�P]�3y���b]�i���<�|=��S��@�s��:\�ȘA�4w�P�uw��@�cJ����sZ$=�N'���L	���{va<Z��Uj0��{:������DYA�Ph��>�#�fn�� ����MN���j�؃��1��� k��dY�R`|GaI�@����!���&}%}�N�K��G���^hu�\�F��gt����U�}����md����)"s��t���-��wA�����Z��>��b��H��_��$�,)fY�-o��,yJ�i{i p�y�Cܘ��^*����4�:Y�L[��(K�� `�^��)�Դ��_O���w&7�RQp�b�ĕ�30��'��rXn��}$��&�77T�R�}�4��/'�G��-��k<{�KΈ�>��[���M�S�����-K��1㋊)��rӍ+m���wﾾ.��I��+����sx?��`᝾�o��y����o+"���$S�i,�Ⱥ1�8�b�Z�Yc��� zΣ:b��1~Y߀k�%�?P�Բ���@�k���Za.R|Q�	�Ǭ��ޕ��HD�p�ӝ���g�� ���i��|��A m �ʵ[_*�9*+�{�`��t�����o-�
j訄�@�B�ּ:���"f~��F@T���yU#�.[�`�ɖ2�����'n�(�T��f��ݦ+M3��^��l�% +�Vp��_ֳ�׋L�C�^Q�7�:�8���n��-F�z���)Ѵ�~��\p�3�����q�ڣ �	[�֝��8C�qf�Iޖ$�Y�[+����Q����k�sV���ܾ�癙�kLȉ�X;�>�<�iCy�����r�g.�
YC��{6 CN��t3�`#GC��Ne��L�F���מ�F���u�R��Tc	���J����v�}a��yQ�^�p$�&���1ʞ�F�z���Wd�MRۄo��U��mz:ƾ�s�r�/
�oҘs��:ݳ|�6�,����*$c����e;�������^���B6�Y#���,�]�c�+/��)^w�S�V�e�8c
�E瀗�'$X���A ��"��&H����x�u��I�0����X�Bbi�����δ�NX��uR�B&pMY�n��@>�k�a��(�\�c�UN�\��s��9�BL�2=xj�9-�xY�e���(����g-���$��:E�҂_�;M��6|+��u$�Y3U=�Ռ��1��Q��t,�@3"�Jd�}�;<��%���^���p���2+��Ўw�/��/l�أe� $͉��	��4�?���/���K1�B���Y������"(3��Լ����.�?��) +~�fj����$^,7���|<&;bb�J�����'[�T�	{�t�P���X��e"N���.������5/�6��t���<��.U�\D���,|�!?JY�_U�]�7?Q��C��+�F�OR9��!�L�C���LD�VN=*��R�h�~���g4�J&"�u��j�M�!����+��q3�r�� b`��Ɂb��q�0e|N6��5�ٚ�%^�
��ٮɌ���$�1��C�V�ܒ�I�O�kw��� �/�:F}l\�2�9J0C'R�㦜�́���çvZ�ƴ�᩿����A���^���_}�� 桡mH��X�i9���f��]�YW�[�t�#��5�jf�.���f�;�h??@,&��Lz��F��29��r�Tۉ�o�%�T$1��L����J���7�����-�2
�2��K�`o8��C
�'���}O��(����[A���ڛ��ԯ4���?�d�����Z3J�s[0i�^���6�H�i��7_���q��d�j�Z I�h����-:ߡ`�:�V��%a��kzYL6��F֐B����la^wݼ���o90eH�� C�����:����M�&��O�#7�6���e�-x�e�9w�w�xIU�T��t��1ԁ�֦�IBA�L1�2,ɺ�d�35��e�h���[f�)��Ze�z��R�jĀ����ҊţZ���3, �?1<��?o�* �J��ʀO'��r�q�xܓ;2�VkyY�Y�� �Ϊ-���ݗ�#���,���q��׾�G,n�y�m�҆2HR9���s>C��i����O�	N�]�S�>�PbK�Qj�7�$3*���1'#�=*�|-�R"����#����SS��/�� ��ܗ}���Y�yA�����FF�1 8*�j��+�jˁ��)��̀^��˄VM[Qy4[�2�����*�2ʟ�K��r
HYq����~��� ����=�E]�"�vD3���LCw�
��
'yG�J'���z�`�6|�AG	�r:Ȕ�`��^/4;H�F����X +'�(̀��u�>�;�
X�KtR����ӎ�2޲����������}���Pm�hw �������,d:r�s|=4�"
9�L �9D�)���v���ݎ>�S̸%'�i�h��!l�N)����I���A�G�R��ƷΎ �x���N���󊒍��O;HZ�,h^�ͫ����!MB�t�X������u����BT�۝��X����p��r�Ѵ�(������C�Q�6'�4W�k�t�ЍǨ�p��Zsuѕ��ݤ�Hx�0��]y�#��C�?��-�Ē�Ř�TX�;�░5C�^�������$^���9���KnC�mRx��`�0�2>�����x▔�l%ߴ܁MR��:#[���4���Kr\,��*ϖ�1��pz�e�l-h��W�ur�����A�N�Z6wg������	& M����A4��>wO�� �l�bܽԉ���q�� ʚ�Yy�_�}VI���{qY���#N{+��z	3 �HVyx|T*7k*��2��Xg�@�i5|�[-;��u	�3����@�ͣ|��"�hҟ:jR�YyFl�z��^u�0t3�Ao�"F��{1J�P�,2 B�8�)�^����+V}�~�x%^��~�o�嗙�!~��+ �=�2����h�W.�+�j�e{��v���� �k�����98�?")��E��Y���h02pA�X�PAA����.��n�СwDI��k�2��~ ��0����SMȧ�j�`�8���Tӹ�*�Ӂ}*A�B�u���N����y9ӿU���5�:�y�``wo�VߌX�O8����� ��*Wp�{����
�W�Y��j5R/񤑁��-������ӫvpx�UkkQUn$�Ta�S��L�my�@2����(�=����)p���G"TU���39�v�v�/�j/wt���T#v*�Ɖ��fr8-������Fa��Z�(X�C2�:8��8��	 p���ʾN#���v]45TnLmjY��/�X��$rV�DT|N�����=�L�3�Im@����Dz�'N1��<J���4@��,C�'���k9��ܢw��I����u���������H�0k.��_Z�?������.�C�	FIg3���£��7e�e6�Oqrt\~�CC��jFɢo�V�F�������?�O��Gq��z�R�l�D�Ϙ��j�I��d��l <)>����8ޮR�$4H"�hdP�=2��g�W8���af3�hH~��l�����gDUzJ���䢁�3��4_;hl���chh�D9� �U)�:@;$tO��K�%�?� �Ȑi�'�{�k}U�o��{ף�I�"wd"
yxb�p}�hׇ5��|1�|���ҶkI�?}ӝ��8׿Zc�-��o��PN4����PEʅX��eg�0�h�Q���$3�'��Db���T׏P:��	p���ߏ�?D�l>�<���@SЁ�o ]���F��F��n��?�A�'KV���!ä�y�b�G�t}Emm���&�:6��gRi��Y��_��[�o#9&$��/��Z�RȘ�I�e`�vǇ`]�(��ȭ]����)JS�rz�G�?|���c3q@�&���ݵ�2��RI��u�Lk.�]����$�cd#��e�&���==On���|G���0�o�`����p5�w������$\#\�[���3-���ZN,>���Y�Ao�G!~�Mo�^?��][!�f�+]��$�Sj*�Q����gv���|oNƮ��>Ղ�x�&b]�A��Yl��ј�ګ}�U�h������Ң�I����&z���v�i�þ�G��\R��\p��8��5r.7K!��=t�G0���$-�}��u'D������S�p{����6��@�~�����ZQ��Ί�;�������q���Kl�2���UMg)��&��,�h�O����V䉨� ��O�GF�P7����	n��o]�=R��k����"����fg|�"\��g���3�'n���A���}���{�"W��Q�2@�:�#ګ�o�8�������?�T&�$%�S�'���Y�齬*7,���yq�5"4~���Yҫ���	x.��!�t'�o����Oz�,��1Ɓ�G�����9̩�T��:�7��l2'��)�''fNo������X��W5?}'%y�7��_�K�X������~�"�����i�$�����&I� W$�#�Ȋc�a��]�Z}�6}�g��R3�s�#m���&�L��s.>��>Mr���ݶ��7 ��<]X�A�i�1����Ca���b��L �q5!e� �[4}�K@��sp��"�8/�#��n`5�P�2�0�x`W;ա��ο�]����hLp�n٥��)�*Ͻ@/�P
�9�1����(%��q�x��e�eg�i�Mg
N���w�
t����| N,h�Y߼&�{Q����_2--�--k���4�m�'b<2�����b���B���^��)g$�N��ؗ;@ ���ljb�Py�aaz��f'
Q1����30�wI�hQ,�$��ω�h�V`?W�],�e�4^{t�;Rưj�(�qc<ʳ�����	��e�
'��Vo^ޘ��ؼ\6D$A��44�׵���u�EG�y٧���O�j���iz��In�i����E^��0�F�2l8�my��垰�B{�,�mq�����ЗN�6�� �O�K3� �t҈����Լ�(�o*ۘ��3���XxaoSd�,|r/��&-���yK�%�OAw����M�Aq�UB�c�X�ĭl�ixh4}D�~(����q�� ��_>(Q��X|��TWƔ�����$@�Q;�WX�wq�c�1�/0����C�/a�u�\��Q���]�j����zs�Lo��z�Ch�a���a� �X�\�PS[��h�?{J��t�[�/"���I��.����s/��zz��9 �ҾJ2&G�RQ	���{��5�$s�ɱ1-؎f��閌e	�X�#�����O; j��i�}����NT'��'��	E�F���?���*&����Ȝ ���<0Q�������c�S"S�aM��(F��Z��Bm��ۼ�g�F!FS�F~j8�FCvnX��( V%pߥNP����%p�aB������Q�����ۇ�t�ː_ē'r0�O��7�٘��q3�c����T� "��p��h��w�q�
^�}ׯqq��\��9�q���]�Zޤ�u4��u�\,��ʍ��]�2�����,:zg4�0p��Υ�{�����=ι��H� ��m0�ͽ���<E���+����#�z��1��^���_�ʹ��/o�їtQ&�L&)��ۜ�_q�~��S��O��P�`���$�p�R�ҥ��n<&
�����������(5��I�U�BT]c E��g��b�
#B���%�GЯ`�1��f�|3��oa3���؇fsm�b��޵��^�IQ�Ah�zg�*�L%s�s:-������݀��f�_�wc���L�Yd��r@pu��JV�B �����c�v�2�������g�;�*W�<��uV�Wά�\�G�@�>*�C $��H~F����m�#G����|�4foK���T���+��i�.~܏o�˰K�#��Y���4B�@�{.�L
E���m�����?M�S`�"Q���lU(���0.S5�Ì�`�� WL1����E�c� ��V����J�N��n��%�M�r����;D����>���_ⵛ�EN��xb�Cm��e����uv+��<y��(m���%���bF��5"�mX����_�}D�_g�׸I��v
�#[&�����-��E��m���ܭ�S��7ـB�*C}V�j�����B��y �����09^v*x4��KK����������B�^Go�bsn�7 � ��*��b30)o�K�����ۣ ݾ�Qҵ�6��f�|Q�Y l=�zv��1���͝���%~�G��#�1b� e�&[Q�C1�y� �=iY��N�wY�T���Du�l����v�<�F�q�M���>f�����Ug�v%��%SdY\��� ��#��> ��DQ��޽�ѤeW]ɦ�ǘhp[�L<4A��M�:�奮��i��@iJ�O.,�L���XE�W����m�1���R��S���PH﹉-�p���9|i�pT!t>2�Zo��Q���c����v����Jm{.5�K�A6�.r_*U�ߵuF0�}�K�dq���M9����WhG6"|����[�]�8�wӠx�!v���oR�YN`c��:�=�0�Nq���Vk[M�=Ԋ��f�Pt_���㍕��<����p��*?�I7�0nT��q��#�-���o9������lѡ�X~�~���NY�����ї�Q��@��㠯%�(w�h�W�ӱ� ���r��f��t��ɭ�`<�3K w���&�Ũ�@�
�Y ��nO1;q75���*gYP����D`kX>��#�����v�r���IZ`>��8WW���D��ѱ���+�[��	�cW���6V��E밸��޷������Ssb�q}�(}"BL)GrdfJ�Ӵ��*Ei_�Q�`�������tOFzud�Y��O�0�š�}gഡ@X��q,s���M.������K&�,qVA��^G�[�Xu�O=k|T���B���x�|x��)v�wӟ�p�+#:+�IS���5Ħ��<oYqV�����&mP��~��H��@��W�`ܼM���ɿ�&�G2�-��o���^��DK�,_[z)}�:�B�]��F��w뜯c�DOz�tSt���ҙ�|���x�+v��|	%��'�t�w�P�閟&'����?���p�@2�/չ��'��j�㗏$岚�]�V�[�ž��n+-z.���J�����A<���҃�&��oP�
k��֡��{.V�h~�)�9�^���U�]�C���ݑ�GY���$J�cn
���r���2Vh�h!���q��&�]0�[��܉�R����䩎x�� �%2_� o����l`�j�E�/'��-�V�IZ>#�6�~!
����H�k��&'�`�V+����"���M�����S�� �i~[L����?�|��Kr�ۢbM-��X�&�-,��h�/��oj;B�l�}(�y��Z��R�_%�o�$}����v4)�^ɿy�"��+t��j�R���tc��s�<ϸZ�k����地YhC���\׀��E��>Q�)Mu`i����"RfW�!q��o�^������2��`�M����9�1۔a��*�c>:P��	K8O�zW���5"�����f]o��^�1���x-�'�<ݽ��ipJ�pYB��LP0��o�m8�����ƽ��t�	Kq��w-5S�˜�d�/C>Ҕf˦����r�8�t�����~�����0�g?�zc�� Wj=L!��6�})�vF�בR�I�]���.����N���ʿ�x��"w��p^��B(�F?"�Rk�*KD_l�^���%A�|.݇C��Į�^=�Gr�DAd-���/�D�j�-�^ef���x<�Ӛ�Q	���u2
�����h����0�(��{���Y��)t�`\�a]|+
]+�_]��R�C+�,x���tR�1������i�����i,�zn���THEJ_I�+H_��~��� �G���Pq���.�C��VJM�co�-*p[۪[�p�g�7�"�����I��<lOs��iI�g����sͣ� �s�,������=�־�z^)#��w�gcY|��n#1ժ�z�F�jpGy�����&1+���S��1^2���zy���ś���JƒY����}E��<����:�<������qj|z�����9��:�7�5���nW�䀹�#6r����[����	A �v�c�{�6����#��59�H���J_%_�C�Bkg� ���
�A*�t��Z�M���dO�7�Q07���#��g;C]Xh'/A�kg\�'ݓ44@��������9�XQ2,m�|���ZT��VAI%*��ڭ#�ф ? ���HK}=���n��ʦ��ӹm���� R�ڲ��Sh����Sن'q����e�j�O��z�c��q��[[��!��ey������,�o�.P����z�~�<�s�u���%:���*�B�r��I��-)x.��v!J�&I0���.�p����������R���%��'��ҫ��c$�h��qa��oe��~c\�i�,�=��ʆ���LƲ��b������a_��ㆷyd��i%�o���	Zu}�f=mVf�8��~�/��u���C�����u�'*�jS��j�

��	Ѿ=��%���{I�P?F��R�w�i��i���N]D�!b"oC4�!]���u���~i���P���N��_��篅B2��/��ڝqT����=b�	��d�����d�'�Å&(7�L�}��-7&��A3]	|��>�W��-���İ7wX�۱4-̎,���ݷ��C���;���w��Ϯ���Y�3����=]�ω�,�r�CDS,t���埨��F�*º jk��N�m%��ˡtv6���T����KtqU+KU'���w��ί(S~��E'n���������Fͤ����Ì�G��|�0�D��)?���-����l��F�m����̯p�f���3�����ى�,��:���
�<ǾVI�j�sG�H�����v�k�S|�R#0��h����k��\"�����ۖ/kõ� 9���Wz?�����%q\��2|������u<�֓����u����}F��YG��q���P>Ž���3��C�����w��ZL��Xg��ۂv�7d��-x��N�̛��"�&�Ka�Tq֕�>��?�.��ږ{�t�;JA}.�N$��u�㱔��z<�v�N*�'�lkG�޹�O0��/j��z��t�BUO���]X�f�6�5׹(jվw�t��0��(��dՙ �~��*����'�`�T%���f ��υB���ٔXx/�?���<�����ts:�0Nt3t�++�c��y@�uڔ�2�N@s�p�q�C�b,y�m��5S,.���f����~-�:��~�;⹘���� �<%��4���a�5�?�`���hZ��C���b@j��³�u���ܙ��@c���M���Α��� ��R�j����C����1��g1{!���QF���͛�ţ�����e��35�l�K'����k��<���X�ЋFG�7�ޡ��K�6��4P>�^�Bb�>���*�,����9u�:�F��ۓx1(&��\��;�4��;��
���?v��*�uϷ�iVP�>�u���b��揂i�X���H�� ���w[Jl�;{��w�*�N��+P��N�^��R;/p���vk�i�L 5*�M�\�c�GQ��.p��YLku�X�:h���D���΢�M�����p���%�v*ժPG%)t�z�&8[� ���U�b/X����R����`_cɧ����ɦ����&���<G}��U!8N���l������tҁz�ј��[���������|����b����C2,C��NQs��9b.�^����@:v�o�c��:��s\S5E��^��"���͛h��-�n
�d�[!�G�I(��I�1A�"B���Z=�곪�$�gr��5A�����dT�o���N���k��4�s�O�с��kCi��2�QĞ�	�#�|o?hz�V��&G���X	�ms��1�~�HT����ApZh���r����l��x<2���,Y��K�z<��}Mh�r�K!H��
�F��xh��۽Z;b������E�ަ�:mD�[�v�"�>*%ܰ6T���Y;ұ��/��^>:�N3��d)-�&����3zfz���MJ+�\S���ZO�>~	\�������Tٕ*<�<�z�'�rE� $��u3sW�mT/��Q��.͎!��צ���Z��b�
��,��g����e�E9�Da��N¢d2R[�Hv3�eC�lآ��� !���o	��R8�2q�k%�О��۝.�1�؀���P�А$ۜǖnzbȾ��N	OVE_�9����i'���XH3����� �d�<�k��JΜe-b�UB�w��J]H)��d�7��Hf�+�UO:(?u'��T�r�`h�ρ��������h|��7�s8pϓ�*P&�R3AJ��`�࠷Ћ���2��H���_9~5'�U���EE/�5Mx{��|�XJ���=;�� bK�f����-�^�[����J��C���n�"�f���uR۽H��c���Fj/�h���%��T�9�/N��^�:�du,���}������\�)�Cŝ�j3�-^��(�Co���i(2b�ȝu�(t[���a3�n�)���RqJ�(�EQ5ga�}���T'F�F���$;}$XG����]!�_ì��dH��D˺��_�C��?K@0���p-LWԡH7��@��v�	����n��Vg�X�R�"D�ڼ�)�[t�rŨ���2;k[8�;�F]�S��������f�C��u�u�I�3dZ	�X�I����$�8FHx]�cNd3he��w�`eVX<�2Z�ӌ� �1�i�q�[���jnNB>y>ƺ:�A� � \�B�ΐ(���%@4+D��V�t*�2��m���	�ފa&B;�ۡ��WkZ�s�7�	P��jL.���~my���?�$K�wi�뫘*?�dsVt%ll7��	���$'���BQ�e�� TI�b��Ù����~����������-M���]��V��3�ΰ\���H���g�j���cPN���%84�����ή�����hx]�+y�����*'i��M�z�^���\a��^��E���B�δm[2*�uA�Kj=�]X��sLa���@�ؿ��*p�iQ}���U�����kw@Mp~��L�d󗹙!���PpLI�	�<�����-�V��c����@���ɜj�Y0'�f�!\"z�w�Y��¤7�d�"$kxy���V���"�������e��8T�I��)�l��),s/ͤ�Չ��B��$ۓ8!E� q;����>���뤭XP+_����IkC�nS���i�a/&��`�C�L� k��$p�t�5�`�F�κH[H
�9C�s�
W��D/ƫ�иj��ǌ��	Y��+R��R����hPd�g���Q%� ��;z:�=�q�_wE���C�E����0���p͘���H);s���_Py��#v��oڍ�Ǣ���K eQ$V��zu��R��R���:�܁X���ߤ^C��zH��X(_l\>�o\b�W�<��0��v�g�]a�y���WR���
��#R�����j�Oa��cp^D�(3�[0�Z���?jE�`�Pu��	�9�W�|���I<QJB����V�K���3@+�8	�2�.��"�TE��L�CT�%�ª3��;���@��u,L/��\9��@��l�O�6a���v�d5qs��K	��'+3g�&�y(9�\mUڹv�M	��p��81����7ԏT��	��q�V��-7,����׵٬���6E�mߢl�ZA��b`�r��|��ɧ�u�����w5�gބI�	�c�kn!s��@�y��K�vs��o���z�ӓ�0��'3�$�)'e
��!w۝�1��ð3��筃��$t�^��<�z�+hӷ=�_tJ��䠇Đ�}�t��}:��2e7,M��bf֥Ѣ+���H6LY,�ֶ�������Ě��$�G��>p�-���Tҫ%�� c��=���0���l�Pv�$G_��sn�S:�SoF��%��?�8p���xI<2R �?���8��VJ�Z�e��5�!?T|=5�M�F��C`�J�'�1,�ھx��<	�`�8��_~EcǳT=�K�Ֆ�O��xW�Ϸ�3V_�u��K���A�&R`��]j�鰰���WW�pb�y�a i
�V����nz2�df�t��Xμ�p>i�_�Wsـ�4�i	iky<�I��I���J1R<�Z�Zr�!u4��� ������	kY�
�g�6\��T�LiC��W��uW֨�v�0| [���~�+�m��NH��Q���s�7�G�;��Q�T��F��H�/?{kA��M��o0�X��9g��,M�����������*�)����Y7��Y��=7��m�_?R��@ 8��5 ݻ��!j�2�?,�e���dZv���^�bv�j��?��a�$f����T�����/v[�F�=o�dP;R�%�?L�L|v}�u�,��V���r��%��o����9#r�m�~h�̮���^��_��SX�p(��'"ų�12�8}jK��A{��������,�Z�E4Ľ��!y�H�� �WT��M��Q��|���w
�:#�J;#�����F}ur��3�+}�͙��x���@�>��z��Ӣ�d2H�$F���t^�n�4_�h��NQo��G��lc?�J���HGC�M>�܁�Am��0k���VK�d�+Np�[&1��Os�>��#/
�\y�M��C0�ߘ1+�#��E��~Q�]��r�^��.�\���2j{�/���&4��ֽ����<����w`��������֛�=��h�><���fM��b+���´)q!*��Lc��25�!��b�DA���&���ƥ�X�X&� �	�_LTA�~Iu	��/＆
̷�u=yݫ��H��֤�	����`|a���m�A�[lo�0	�S�?�R�	�i�<��e��
*Dk�����)�q��'xÕYd�`sݒ:1��Ѷ�u����-�NWM(�%N&IM�gr\Q��G�p�:��O�ˊ >0i�/q4���+5�:�x��^ɬ�����)O1�Y��=�}���fv�{����p�"20)f�b�R�!S+1#�ep�b@VPD&�H�="���ws���=::@uH)^H�bw��2i�[�����Or�	���'bd���c���P*v'3�w�\*�P�J�'&�Wr��*J�����#|�!8�y3�{4�!-�GBy��sj{�@ Y�q�
�qO����'�6	�I�:P2k�=�g=]x���!�g��.���A��5�l|w!��m8���]��dݡ�w?D.����[�����vZ��
�����ϦgS=����,���?Ō��-�R�Wcc�[RXŰkM����;h�Hvv�7��=쇓��ceu��A�^�,t�Ť�e�|j��(�'�O�8ߩ'�q1P�j{5BSh:�zd���5�(�j������i��gѵm�C�(P��Օy�$<�
�f�_q���P {K�ș�3���fa�7Yhiq�|�&[�V�����@��Ъ�E��O�������u�)DX��-�y�Z���>١ �?��o���#.��`�U����	��bK��~�e���Wéݻ]{Pib�`�zs�lP��Z��<[�@S�8���:~q���)�$�c%�ң������5���k%��Y�T%��2Sj?VH������@�&u���ș���Dj����?��Eb�pml��Ŝk޻~@1/@63����(�!����4)�������U&>\��\a<���(!#pE�S������Þ�JS��E��yȒ�	��.1k�I7i��	�%��l�Nֺ��B��3Kg�Zq�&���>ʾ�;�m
8k�3a#�]�0���>]o���bn�,7O=Q��r���DR1�g
��͕�|��Bu�Jj>�X�Ls  P�*TPf�(�N���)7��)4/��b��� !k�'���C~� �!�����E��3z�Y�3�ޕ��n�e���H�+"Ex궃����S.������P+!`�C x	^y(�&[�(d��e�b*B d���� �z���s�)�*���;	W�Kc� ��F>��'�����Ǘ��4���}ʆ\��q��]����[�I"
����M�(g�j���5q�f?��kG�)� z&UĪ��ߕ����}�#��R=�����/�k�V�pqW-i>��K7A�n(���]���u����q� m�lV(ٸ��#��\���d�Ŧ�(��g5��s�.bxd_�JT�>��&��u�፧�l�x7!�{աKJ�I_bN��Z�v���E�B��ϙ���V�����z���_�a�r9���/��r��(7��O�L�J�u�N���ȗ2�>Xf�OC�ۂy6S̈� ��V'#3�� ߯�U"���n��)���&��K�4~��t;"�X�Ǜ��砝�W��1-ͪ�7�l�]6��V��,�T٧���M�lY�@�֟��P$F���uXΦ_�	��Ȥn.=�v�D��m~:��r��/��};ab�(�hk���K���9��H6���u����<�Ń���JVX�$F�f�15�y�A��u��pi�z�RՂ��<�|��ʴ�C�;���GH�[�����5�u�U��/\D���ʬo{����VB�Q`������"����^�SI����Q}�QM��k\����	e�'A�aM��Nj�9���Q����;@�K�T�*�5s8NC�3�/�Ź���R59@�IM1Ó,"MUH���;Y5�dtoU%'=���a�m,
�s�rPNm��}��v5D�����t���vԼ����8)2u�!��ʹ�Zr>n�q��r�)����#`d��0rǙ�Lh�J�a�Wgj�p�X�����;"����/*��A��������	�|�Ƀ/b����Q��t�wZ�-�_����}
b����4��(7w��`�cq҆�L��&��v<9��O�r0Y�dK��XLj,�l� ��t;����u:�k�k�p���(
"��a�_�Hnv��a�x?���u\Z���_J{F��)��I/	�1�6���Qo�EA�W^Q1�ٵ��b��������:���	�D�d��Y�����p�~l���rZp�^�õA�r������gE��ڌ�2�X�E)Tɜ^��h�T6[ʹ��q3�	�C���K~Ҷ���e�)��I��X7�7�,>[�����Ifr�@����c��cd�H+�h'L������u9lbؑ�+sˌsy��О�ҽ��(l�HKU].���~Bj�i6�B��QAk~-p%QA%��d�]���Ң�?�׼����fê�i�M���>�eΉW'(�OQuc7��>���S�v�����q?#1r�u��Ox����`�̯�$$�0^��$��̠��[���m���*�qp�ITq�ԤXᙧ�l��y4P�󴕷�wltۀ��泗'f��eM�}���!��bG�7nߡ����cYȃ-�Ј�/�4Pƣ���#Ћ�V�)	��$����36W��V��~nGb0���Sڧ��ګ\����b�t�+�Z+��BO�W�==�$���1p���	��e'g�N�>�d����n;����q0|N5�J�b�{[x�����÷�2ӟR�H���:_�S�9!��ZǏ�{XTjOb
����S��}��M�A*�ar_T[q�Xe4o��(D��y��w��:�F���ㄔB�T�~�m?�/��ȅ���c�j~��0?��DfW�����5|��!K�������0�6�_�S	�E3�����۰1P�.�m�2�C��|Q2?= >�#�B�~�m	\sQ1l�T�L�HQ���C����?I�'CB�m�j��k�/�6��d���R�E�Qئ`ݮYB�
N�c��IJ���k�M�a?����eX�3V�ǨꧺUm`����i�|�zg��@HR�]<�JN`��q��W2m����X<b��F��`	���u�QH$g(��a����IsN4)�!T{cA���7ԗ���� &tI�}>-�@�^c���M0��~��_��N,��s(��B�L^*	>�3{���IK�0y��|P��P�t@:<}o� 9������f���#{U�"�� �2n��t�I|
��ؑ4s[2�����C�o�e2���w�=�<W���h��>5_�iAװP����(�#��/��v�w���Ԝ+[�]��d�ү�.߭iKa���%^�rb/�W�T�j���[r�����^.E����]ꞥ���2,��v��D��,h�/����9�=���NִO>?1��� �J����#U����{|�)���{K�	a�t��+�M��*���� ��W(�X�0��VX�J��R��GM_O�ѱ����A��F�ҵp�����ْ�Ȥ�ޙ�ۈz,_�0ߓ�a ���0��DT��(l��-�@�]R�mB}���$��r(��o�<?P�	�/���Y��So�}pt5˧}*��������(BeW=6��D��-'h�����/��o��PT����<+>�ʚ�.F�����������S�خ����1��I���x^J��A�i�"��}���1qdF���7�U����bp����Ņ��w�́����`���������{�潽-w���e�wR�K�,#�Ue= �����!Լݼ���T�Y�[U�S��~|f�����чM9VI�V7����������%�� ���W���UN	h�u�fj�*�0�����P��E��pF�;6z$Jf�9	X���Br_`�}����Ve�YCHydT,jns�u�r4�m��0�ZgU���E�:
�����<���8���!P�Ub9��sP��ݤ/�~�F.���J�f�6t�y~�r`�:��ŭ#�R�Rv�~�H�rL������?�z�mE���P�a�	
-����8s�]����Tq5���Ǹ�[F�H��~+��'{���	�Zv.^�����Xlc_e�2B�b�>�s.yoL�'@�C��ҍ��("��=�WEo���%���� ��}�ٴ��f�G�([���cxɣz@���S1x���m(�ᒚi�a�!f�~-��'��X^9�?��PF�{��}�
t�-}�hpp5+A
{V���J��jR�xia��(C�`�,jJ���uu�kր
_� N����uH��i����+VJ�K��F`9(0fm"=�i�����'j�7{��F�j�H~`J�^4�vڽw�{�p��Go%]�x�mT�QPv��I�(tЉ2�"�7����eOѠ�`<�C���e����������YP��u��d���x�~��%5��.Gu����QGR�3_Iz+<R�"�� z�?����d�y��^����l�LNd���ڂ�+�i���xu�䏋+��[le��a��&�Ŝm[�{q�p