-- (C) 2001-2018 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 18.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
12BxDXjLY1BU3JfXnCc/7GWH/IGBc5Sg0rRMc3RMqxCZMh20HlkKtYsfhcCrL+jQ7uA9Ci5MLyTD
2OveW3Az4ZdGPdWuBCfIobkfY0sI7zRTm95o7PSAfKgfy6ZLmiUqB5BD7sR+Dc/YQuXlu1E2qQNR
4zLOJYcdUt35gHctgmZpZN6lP/a2zjXuZZK6uPmj3pkwSmQwfoGCSXCfjvnKzW1OIz80IW92MH2c
KmcqDilIYxt29Md37eWoC0iWYPa2f6R8FcSmgKmzkKs9LvwjISZGINnmxPNQAy/09BoZqZB5xMqb
6UsGAASjPiDYhI4RMbXY+fDHKRE1gltBBWtZMA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 17536)
`protect data_block
/zhWG8OeIr/TUaQqCmKAKDv6OpcMaTM9AOuZrIVOOhf5aCiIhRDs8bwOIpGLcVyCg6EM0u7cUS08
GTbKx1Fc3tu9B0XBcyewTN1h4eVgba5xd/oubg70WRHMen+RYuCoLPUXDu/2+sh6pTEwiKaDHUKi
G3T2TyaN1CYhvZS+DBYaCUIwztKvHCJY4G/RdjaRJ08NwtQBCILZmn4W98l4ZJRxyEoVZG0UVYEw
CG5oqwrx4zlY2PjCnda0sLaezdr2EQ2Wa82JNNAloDpJ4SZpNQY3qVtSEquZD0Yz/e7SkVccMjIJ
IVdE6x/duW1mX+v1xUxzIe5Cu2TvEpFLuHgxVEmTGwbBxgzyOETSsex3Q35Y7gZ7Uw66QQaPCgbp
8L6RmBIS/J3/4dttPc8b4ERFX5mlUfElDg7X7sFmwzkdEBldisTbVYdDKwrXqb//g2E9hqcssTRV
CcEiWgunZ0I1e5ocw289pamD4OZOSRlakIrip4mSmhFKlJa/B6NTW1XLaUoQIpxfrYBnaz+ZHlX4
bknZ4CjTXq6uZdk77DUKTVjuPqIjfKrvfrEwiQRZrSTd5PyS9TCWxlyq3D3ei0j9Gk3LQaxxVL28
AcPndOFoLh/gYdmtyqh0EK/37oIPJ8V/hZ7tByncZxgKUR61BWQTGI11Cn2ONofWoY+3Bn/OcAj3
HGyQBUdPnQytsVelNF/dbS9/xL+3REPIQ6tFoLuEeyCC4Wx5+4qSa5Mpu+Xx6Zl2eWfzi4Iv4mg3
WFm/Fh5q2D7rxt5jHoksmYzl7Wq2nD4xwQ32PGbxcoD2dauZ50uIbFX7xcBRlx2iGfGcbxVhGcDf
q10hbK6NBzb3Cet4f4yKBmdcAdFgz8Fm8mkU5m09ocYfrvoq/2eELN4sl87GGrDscLXmMha/QL2I
8y0EFb9eQYP3dOxEZgk/+jL5MLF1adWWbWnvbb8FyXXMI3fJVIkA8Q3U+djaNeT4/8G0jiTUyaiP
VBS1X9NbM5+njfv/Xrlh6JmFYZ6Gp6ptQ5f+mMkxAViTfeLERJ5G73VA67JvbdjR1OhHtmUv7n0E
NnG//9XJ8G2/JO+blDLIGciHhl/CnDtsPLekUOEVC+EVXY3fQVaFYFpq2StWXbHbXdOQbxrsCSSX
zjxKeYmYQVU87wLdPwCjFY1vAQlqlk2lNswBjOoZ0gj6CJ8QWhFg85BfoFmTHH8D/gJx1B1AMYut
mBPYysi9vI5VdUsuiBnyeMGSz7Nh5Gu2qVU/z9HetOEw064aUGJ6LBi7blGXKtyqixIna77nu+IQ
zMbmSZ9F1scUqMv3cOia/ULp87roV3pxReQMpa7qZKSp2O5mbPeVZtVHpJVAYK68Uq7YVqLp4BEu
zu/IZwcG2/ImOayoqTJc6A7YrNGmgw0UTXLWGDCqjD3+72LsB9CRn8DX00M/ixH0qqSAJIdRfjov
DTqQkPbvCY2+Com4JmXBIDfqpgM7umBQKPzD3g1PXQBlIJhcUQatnxLtz6CM8+V4+gKgL4mu+k2l
Wg2NkW7SIdyJvVpaKqm2xnijDzn7lwlWX9Sf745fOWDMLWLm5yN/2ZfAPj9Xw5pZ+2ED8ilC2vx3
oUzctpEfTqm0FquD9asw9qpbeVs1RgDshFkI9ZrENNqnob+xMScOqqvrpasWKrw4HqJG1DEAzfb7
35jcbkXBFHiqTxUNqCUiVqk2HuLnOtIwhxHNDXAi1KGF0aQ1Iz5UgTLoGQVgFXLSLBq19ejGMRda
YWlZ1L9GOZFU1Kf3qAi3wqF+lIV0Qjpb+K0BeErJw+rRQeWp29Srd2KhmWIYtbx3Se4n+wMMjZtn
qibm382UXtV9e3WGdDZyGupDH67EqVYZNe1v8mSz5qWLj49i7eOnGE5N881nEQI9R8CqNU3znbkq
TuhAJnpvW0VN3CTfZbeFFpJ5DzPZbVcabAEWE62DA4mgcZHWic2+KjkGr1ruJNPFxhuzUK0MFq66
QsFBZ10kdxVpJDvO7QkmmcKl3vaSF1KQRFhxdRFo66CfyC9+Dm5RJkyakNW8lKGPPQZ6mjkgZ7v9
F0MBE6cszpHBSEW2BkRhIfiliuD3p5f6/ShwgTDfjaRVjoJ7YBDNmD7XWKRMu0XdQpR/KngUjq/S
NIZPEjoOa8kp+RlY7BreXQSfP7e5XMZdMFa+StaSTo8oUDaH9DNunDwx3v+dTdeP64/NQFzwUo+d
NWjsvBlFCJDamDo7EAKOeSTAVCcA9RDUhq4h8NqWaS4D/JUU+BKvdInvj9FDNS5N0mQVPOFdzBk+
s7NGo4Ja5PaK3/DwbHb1SrQIyRt9eVOyaf9lAXqZPWnW8y0SFN9PUYNqlZc3Y8r2ALBNa4JzruKX
hdaAly3eWLa7t5QEzPl059LAn44nKgmdig5A0IalVP56XTp7NOb6La7M17qF9l6BXHxysgAexxTf
O8mpHEdFMsDZLu5kkkntJEr9o5zd6d0QLZfU6yyuh+KNR1HUoMXGEmC0ufSTm9OnNPsv8SCKQQBH
I73Lmhr4w8wSB4RZdqBZDr2ZuP6FOxNAhh7fn2x+L1W5I6NpMNMFAC7kDp41r99VX3M6mZgANo6/
0HTSk9J+dxMtL1/F6XNwTxYHoKWSKdfcQXFXIn2jMOEfOPU+R4RAi8BtVgq/nii5vsxhE40MzPhd
aSEgNa6eK0a5n4ErcpO3eMDAvw0rOsdyYiZ1INggrLn0Lel1AGuvx8JDmaoIjh3aGJn9AGOqelFr
0n9EIZK2R79uSy4w0jjjR95M5x9AEKrmD6QIHnCl6dbBbUp+vGe1J6XrbifOlmahXl1oKu8yenF9
JQRlrNru4ybiTHhE2xfyRimzwDsZPam3ol1y5I5ZUAp4/vVjAFcCWxyobfqM8ERlGU9XfyKNo15/
pcEaSC8kYsdgm5zyDVw8D+dBl2u5tV0E25gerATA8Hnqp8/RkmX4n97h6tBVeT+WWzUFBimyJ5P5
lHKeq7Zox+gKqYYFTI72w6lY0aIP6+hzbneDsBf+w21Lu3aGTO4VXtz6Z3wodRMqJoy2iEY4QaN6
5wANMqqrF9mtf1npETMZEwz69Y6gBpmO+qdKTonuIFqwazoUiz1DAwhNI0ZlsMqiLQQpNsCDM3uA
P+rL06YjKSPpNlngUepzsA5wZ0xpmPPrVqwpIOGh+TwBmYocEMDCXxW7gP7dw9BVuxC8B43kpVwK
udfW9z3N/Paq+qAN3P8Qib2dXi4tg0iNSAdW+NiINSZw6n+8IQp7zccf80860t5RXuPZy1bnOz8H
1p12iHcyJTAxASJjxXpWY4M68Mj48jFra7UWFBWfttUO5fkhMf7V6yvbEmGIlRS2QLi4h6WPl7sd
5mqp++Ck7lOkaGpRs253lN3Ki+hdVNmTmdFAjFa32xKphgU5hlT12Cz6A5+isU8GdNS6fCiuJTqu
HoGlwWCEbZKVd7pMLJuhPGKoYldKJB84r7lIirn8U6hRBHHYxiI2oQcNJCVVFnLwKEVNDOwuIbtE
8TU98mJtT1JnR/zbkx0UQFUtPD1FHipj4yuzAbtxIq/K3G1B6gROixB4fCWBQREs/lvg7nfRevxK
dMeyNdhHtAQAj1oz7GcSGu0PXMNQziuzybLTHvJGx00oTzr4giA5I05Nf7H3rCWTRNvWaqli8dMa
/7ohztakY3yKjlo4wD31sG/rm5TV2UkQSkw1F88asQpsxvRuABth5hB+IArwv8QdO5zB/kLvvR6w
nNumkV6CzxK96AK1WOPOn2nsN2J+T1Pgwj+o4fIZdYhVxIz3Mv9dmYYRONdK4NUimIs+M/ycJJiS
sm8ntOJV6cFHOUGT9KLfNdrkzsSIIJZIFi8um4LyK2tyDh73MtABvIBKr0u2+6JLaATI2TQ1rRJJ
oCrNGDMC5iKZE7YfVChQRVJHeRm5WtHAl8gojTmAcJ+kZ5whKQ0Y4VQ1NMjQnn35sUx98+oQeNwd
YvnJYPZ3aB3TnxSvFtrQEXDSjqFLkpwgM/NUwGruTXLH92OmJphTflgq8zJoUTDPqSfKwE+PoOCF
tksvsOHsecaVsJGwknHKH5LuJTxdpC9S1N9thagLgh0bj2LgjSpCOKPprkKRcgsISqZAuNgRgT+L
uGUP1T4NTcydKE4ykw+y72EFhkmRus8HJluYvBigK1Z+ejWtRNF8Ik+BmLue+wMI874/a/yuviXe
XJs1elhV154ztZhUIrTP1VpO3gWcz6Tysxtv3qNYp57r5hQXfaDa4vlr9e0OrGQJLszzLa/1gerr
dOG7D6d5lh13idSt45hHKi//W/61Dx08XDf3yhnbhIbIuYcN05UBmt0Z53nnrCc2G7J5DMyWnKiW
7rtG5S90dAlAiPxnw44o5wMBGsh+N7n0My0hs9bKgKUb7j/Uyq0oMlg4bPOh4AwIqVvivcdQvgrL
WRcJVpc5ccBuSFd5QGgTfkru8oh7IxtxDy23/S2ifoTBVmDFou2SMaGMcQ9ADoKe6fgiDYmIlmyG
E5ap1Y+7SgWlf7cGKtM+u4bDMiEYefjHKKSJJ93sjpjGo461SSks72JtdVwFOilUOM5Sh1HVZacp
oBsNSQYSul8+Hy0CpjL45FkCUhlEW4hlemU5Fb+yvhAxSeMt75ggBHilkj3GJEp0is/Rwztj5iW/
4aRXsigfnBXltV/6QXjsL5DyDWXTqoR4pcNAmynjoBUern3q11rdEPzJcVqbUVRNYPN6YH9bXKuL
UwZ3qaMC3xFr2qHFyrnPUNU9SkneeXhY5TcnBIYlBlWEHBlzUfqIIZQbvmvVani1EgzBUfqaWDvu
B9OcfVgtlEJeAlEToMur3lfN2rg8MjANtUMRYyViw/S0ACFIQnlJMGita/BRSq7+TIAqmRmhyhdJ
SC9xT7n9rRWNO1q3DpCYRZqMAM6qJkWHCDpNWQEjDLnsq4opKbNuvKeKFCEwRPZfFKqBM0xPgMOZ
hrIBP4Q5eYK7khgGw/QOWoOV6tpy2OlKUmvOBo6i9qOy3PWDv/apDAwuMP0OhehyBa4nyUr/4vlw
vZS6QqVzE2rJuYJBVzB+Ad9V+haSNIt46nZfgFXJPEmXhCeeS6wGEPEUmFRuEJ7BYVPHxuuXJyxZ
+vS2nXxRLb66h5CD8pRNSox9FgO2s/TZfFi/ovX76J6DCEDncto7njY17uJ/sf9frgxzjezR9zO9
kUe1wIwEN38w92zvxu8q9eyWDTW0sKAJ/WwNWbFyoT9jN2k+JyZ4xrFdxJbjKTTOIOhcJvKdCf2T
YUqix6UUP7BQGEfdvpyPnDyPPdb9xH7jqATjdBdrtpxaEcKUJ8sQHARmmxxSiySdpB7OZUppxID5
qD6KOV0eCjAD/VJCSJJyQH1ETLvefEOY174/wZoFTH/mPid5FPiYtCoC11ylSFy2xCHyrF3hBQll
jicXWH4BTnvrg2+C/hOmHB067I+yyp/kI7lfRWCVU/Ed0Uq6LQ28hGa67qIUkGtn6OXnyubqGLIB
4+b1QH19Wtgd4JDfPvzmT6vsE2kG7AN9i2p6rLixl5UFpP5uuOqM5rRq+ZIlvlnjiXaAaC9zH6Fw
eyVp6GEKdH47BWPG7r130Cg48ibsB5xggd/rFLk+JwBmShb4Q6k5jV2cA2ml9URXNX76EPIF2+O2
u6Um/7iKkHNYNh5UVwqholNtOAN1lSyp99aN7hAo9/iIY8y706n2dMtMS4iy96bK/B1+lxHmhn9U
77qtp0ZZJBAiCkpczSp9OA6E3R1sHZzV25sQwplrgrpwPg6Oc9p7JH9h1PyJIcrTwCohmunaKj1L
4mN2B7hJgGGkC2lhthPydVi/UiVx5yRlyAfaJx2CR0O0EQTEWoVdsFM8EjxM7R6XQzaLkdpp+os8
AS9vxYUfOkBatwU9O0WzDAUmCYg3N3WolGHJ3+o+YG6UISRDIYpEzXlTJ1Hhrn35pj/RLzcpCUOG
11L3GMFBA+Y7JTZrDeAdnoyiR+IOnaXcz9qk+nrZJCkfzSfyB0BD+IWN0z4wr+r/RTM4KqMiO+cr
i1YpDs91JHirq28eg3at6a6hovbT/0EzL77DD3bgkTTMCgN6Q98TEgqls7HyQcxhz7WXyGwdvuBn
K42sJnEQ0oGLHBrnBVgGQIj10ns7IPf/UEISO/IAISV9I9JBkhIc1iVcbiOryDTxuLDufxto/MN9
nh7928ay+h3PCEkt7jDmVwfVH4oW2FatPigSCdqqqdTjAeu4zwwM8754E6ZQX2cuf867G0VL+ZfA
iwQD41uDbMYrfDW2h9ksVJ5fXdrk5neY4fl/lLP+kdT0EvM7HzIEDa5T10bBEQznYKuO0H7rlAF2
8GK9RCqpL0B/xYfWU+CddozhzPsyVfsGShSHzXv1/yW8ks+TTx8bQzDi9fIIJ1oiHCNHEviR1eF6
vx1+l3zfnYFyemeBQlWIGsY3RFU+LJczgOc5KV6w0Yan/ZEnMqaxfegsOeac/daHmITeDKkLBXMp
dyHzg1ZHJLkuaezMIbx/VwyUkmKDXTKgVay2IhF71pGY5VBzwmjUNihgx64lKv48iJtsRnuaxs8l
0qCHWxlsdFk3iEwoWSVvkNWvUid2jXWnwdz3qwS4hTiVYYcbE/nCcxXt6SGMhmxUBUVK+SLs65wV
fvMdCzpFfXwQbETWi73h3fZOFZ/a0XaFxVxhtAnesunRoJ5vrfP7gQmNupoN1v80VuBHaV7WUrF7
sYYmL4roq5Fu4wNAAcYcgIXPKkm8p9KXkuzSkkQOylsRd+oW0RRL3G2b1pCXfmKWdUhLy13a3xhy
xfgdRAbITwyXD9UdJeD+WdQxefliaevg4R6pb276pETiJdFvBrTLBBZRgBdGv/9QutflbKRk1VQz
n9a6SOAa4ycc8+z9KQZSm1jtIEEJSvBLiXfJsHCX4B4miN2LmwLpTN7yoZmCprKtZwqk+Cxm8GbH
NYcHYJCeXfe9WvB2UfZBTGA+dDGssUMpXiBfhuV2a0hLpgQJbaMPIAjoIG1e8VpBRuV/WCwuDzKH
zg3EDaTLNkLnKrAOojhe/TYBdpzJS/2/PJcE5JG2sXtsbvC2g3HSlFkhbinf+Ni5hRJvfXKo18z5
yz5cBI8JDqQ1xTfakVmUrdpd+LS9Ud2ftu0sgkUHsDYBdhKC5ANDlWSVn9CcJ6BcBRJXblQ6y4wc
+pAIb/rVqZ2OtBkRsyoSmJFpq5wRFR4AnSHkInVvD6ob33x4G2IClg+sb5dxhz6izOf1nJt7Z0oI
CtReUpJzwtPTaNYjdjRJ41EOp5/dqFUgWPn6URi0TRkrGZj2f5bzWlwTLSywKww32j+/P1SHTe2I
QvvTwZO8sMOD59nrTKaDOpyIWEoR/ZXH4B6uckdC0H39asKIArGFZjdI7oSlTuep2DL+BTCA1hj1
c6jE+sMtIXZ06uQRDile+JXQEcMLvmTx5sD9lYfn4iYzPizig7dQchpP6euDLnYKlk56R2XwigM+
20EORMbVdrImEWxa3vGqIT8SxEZRtIEsf8VIfwXpcbl3qcA3iK8djSXT0I1IAkM+GX0J5mDRCoRt
Z9jbYlDTYBi8mVYl1KkniKVvZa1fdnWnG6Pw4eZfdz4ys4+NG/pPO9JHj8JUteo+HqOrlDiO4mbC
gY2YfAnvgy81FVIRNKa29UcOli8rb+/SeMDp2914ZBUfC/NJbAYx68ywTlDof1XRd4JuTIHNj43c
cpyX3dhTuopFUxVCurRIoSuO3/WrkcwCSktJptLcd9yjdKwcGGrp9QTKy5FILZHoQg9iaCbpDkoZ
EYzfhJjfNlcYQrZmuWy2VDJwd8HRGDpOFTjfmPLZ3I5JBPOXK5ADc71BaHJUYFrxv4bkB2rLKmsh
XBwpqnbAlBCzxs0uuCnRUkOgR493OymslyY1I8pLf3eeLwQWrTUdzbHh/jqNok9mSAPuBI3awE7A
c6aL1b7cFhbfsaz3N0UeunIZEd3OnyOf6cLSi7Ih7Rv5tauit3vIKmsplCAmDxZD2AM0mdG/mDcp
RBVXRPD1B/DSKsmDVRWhAd9o6RHSfG3czaRRhDEdp/iBG1q2Ir8FKG4q1eBCuOhZPUPJKGPEDtf0
PN/uZgh52OaHSH/iF9dvzbue84Y+PWylEg0pnQj1kdHVhv5DH11ZWtbtOdEudIWcRvexMz40xH4D
r8HWovlikPMGP1vWwEzlB8ynG/pYLWCDfvtbyiAnsVmpr3BoUigML345JYE5KwVUW24+vZ7rMZ+b
C6j8sBBOPr2IS1n96qrkS7T1HofghJxMo2OhK0Hb/ansnN38WoVwJ3aMrG6YHbrin7zO4o8Yu3O1
Fk5VqqvzVg8jopj9m8bpi44frpPK7L3i19Mt0pPpWIo3qbGla7eJP3N3v4pcSQrLZKRtvGXIJ+hW
QFhdX0C3zfGVZWu0XodEBTrnY6Yvsl7riHs/eskdhQx+jMEhIzaksO7YEchkYEDrGCJI/tPPiFqA
mZ0wGWN7rtme13pqzf1BemUR/BMtZNemQm3+EHxwT/9naJtOvFDvgJlcJ1vN9QpLWdqWnxD7MPJ1
HAe9w9dBSaoo2lF47AFCTphsH48ic7WYoxCbIj5es2rFDQedMGVf9eWSKm1R5wl0oQWhc6DiNkUm
YwN3mpUaGyAZcvQ2GIMLXcY6bSsn6ln1DW9uu+7DjFO2zQSJGwfMZfZ4zCELh5hAkheWI+HXbp8m
GVSooc5rtyDSFY/4b42lHCwspQxlFxURmgiHos8RURBWTP+HJvPA/8SLNlr8tkL2YvIlCv/87vvI
+tTFykaR0PPQLJjEgQPYd0UVbTxUbqTs2sSTr5hMTi4EHujJsTv3OIxNMvlqR4PKgKDA80SisN3k
ZWf7lvv862CExW1WnIPNCzQ7X6al5a3bowhz+4eHXI9rJ/7MC2U9zOHL+lqg47qhtgpox+42oKCW
ohf+dqe7KTU502748eP/gKXOVTeFlAWohQlX4npCXl0RPKWdcaIixht2vo1OMQhZcv29aFNac7yS
F3YR4uUIOHViq6HOsfBi5Lf4umCAwbWG4T/j+cWeGaDRb5YkV1l3kiR/tmxlFQYNOM8LLmD4lfFK
ujdnshowZFKyfGpaHz99noXD+6sEoGXwrnfpcXHwd9Rn+M6XuAuipHjR4KsQiafBMPDyresou3x+
qycgZT/8BGtpAwqcMeh7MkxMSOJMAGQQME0aaFD6tInfCV6ZGeuCR5TKmT9PvZTXXbaBFuuMidN8
4y9091hog669c5r1dlwlz0KkEgg2TNVCyypSYard4q2Clqx2hQcI1UAmeD8boW63Dffk06Z6VBf3
VByKJO+ej/FPg7M3dKbd2H9LU7n4lNB4bURvg/NqMpvZNn9SGkj7bh1moKi7gLmSjNyYFmr5guXE
FuUN+oSTlP3jF8yI1xKJJCfPNUaaP7auEUsUWDWVXiPVB+XNgLrmlkqFQV7fl1MJjiMdyUMjIdtV
V5rmdgauytXUEXGPg4kWcHcCn+KjqUhnXiJYNnyaY3UO1Ntf7KkU5IzC22mn+E1TDqBEDTP+k+Xf
Q5mKsVJzG7K4hlDuWiDkWn0u8Yvmm1ATv4bTI3OHloJSW11sRCS5zI8cTRBsve4ZPJKVtJzZD8Pw
vWdmyj1wH/yeOLIS4GQyy0BPZGJhWbMcHjWBldLugtpOlMfQiFUzQZvLsDdTTcKH8GbSe1+ieAaY
jubEZfXd2hZzzzAvf9lHVlLERvbAplAxXqNtzWdS8Jm7n0UuxRVEC+/awXHI51qvegJDBLB+GuZf
+B/9K/BopVhPvpq+dTtqJxCG4raYavyoWavVtLtsldhu7/a/i11eTzcXRIaQ1RfXJcLv9pjY5meo
0smqqlWd2umYJJ3NgviYO5KBC1Clyli9jySeBZYHJvI3epdCoxIXWwyCLuuyZVhrorYg7y36oEY8
MdUQV+2ccAo8WQh1u1sHEJoEZVKdg0E4for/nYSrlafa0Qbf6mCn1vSt8K59BXGmz+0ODV+QoECn
Kktbkgi1u1jYkWabizmcaoCVQs4kilBIVZI1paT0JkM5OiajVFjLWVb0qxeYMA9ekZtJpLaUPRZl
TVdf33xIyZDiW7R3iGZ8KgEUe/uQRTgKZnLfou8RQ1cadJmKByVVRpB07Uylb8IW0mRxjYZJ9jUh
YPfRGtsSq494p1XJ/Jl5GhQlLdzfNSk7aH+w4XMitXlwDluf7wDMctkbMVOe6UCKek760n4IeG62
vdmz5zRZEJFiZjEy29ILkrzjKxV22BcVIHwenI6TKus5Qf8mlpDOE5VJq/FKTOd/K/2XRq1bU4QP
o75a06eeNllIr0UR3QExi3gWpVQx8f90SX5YSf6T0Gd+j+j1W115cTrvQ0bdLEXZscS2mdjASn20
/37adKDMUfvJvHdRnYoTsCjf2pEgBJqMO+oCQxLJOIKpg1Vrz9k/ROne907PGZcJWS5kvA/DgEGg
Px1a2jeN9K3f8VKZDu8gcJBSEHEweGWVaUyv/k5rUHOzjmzVxBslI+CJQUC20xQxsyy6b374rZUW
LwJeDW2RLEAtCxOgoqtBe96E90WibZIgEDrmtiZpsHnFQ1D41xDfDOawFfPpV1ego45LcrHhelHn
GOLhwkfpusNb8VvpECPfcL7jOPPJ9KdwFKQQwS6uFk5pD/CfcTV4ptkb+1NoZtL9kNLlZn8gSt5Q
zKCqA3Q2Y0Z1vZ1p4RzX4MCPa5OGNw3U8hu3u0jR1U/pcAnRP/V5zUKujJvFJgnwGodtm6pG2hn/
b1WQqLMJYS+JlAZwdUWS29HX8uhoK+07IHAig9HB6ZOKHWUzh1Pf7Pq701lsFRrVosTuz004UCmi
3HqOfQPUCWIvZFcdBbqJzywEv6Nk8pbYD4TbGU4DYsT9QfIN3ECQKVeJidZbzrLwBi/H+d/v+xWE
Pi1Ud45GHCR/ezzd72kjPOjKPnZ0XdI+n0xuRbLuet+T2OE85fVjuX5bUD01FU5/KYL8cSuA1wkS
BdI0wNfQWdn9MMrjCwBCR07m89xc92fU+1D6DM7j7UgnSyf7i8KM57t3taJlGr3h45GAu0WW18GL
5ZHCX422bGzK71gbzysitwvOlmDBYtieVBV+6nN7TYe/yWT6BZb/on2LkaXU73VrS4Jm5JJ7uTES
+n13eVj4E/HGCTnCDfM1uan1YOm+vI7gDPm0GHn1jwQfuD10Xjki95KblIbV94YcOg3ijgHrsGcG
tXmTlO25E+sHWLNO2E3+xMHTF5yYs5bHNLumlArmffa5wEgA5lJ8kFY37uiQk670S9KC/+WGNH30
bjoJMZzZLvr33PqEqW3j/HVqXIb6gGPY55mp7Gs/q34RBb9pqk9JBzCILLhmIsgB1WSO1QovFwSd
7zr7nwTyW990rSBASjsapdxa89LLyALh61rZWnCV23wTuM1dxgfX76dzwmDVehFTsiIT5PEjv8S2
KHV3GQ9tyPzQFfZRz9kMNPkkJYigSOTAFWffVeq4Auk35XG9faOChasJ+Dm7jsHpVfivxp88D7Kh
fFwYyDB5Tp2dGGpT6jNXWg5aytxJ3rpY0cslMthrOsQbjMhlnyMmPlounk7Indvozkidyednlmyo
jVr5cZgSLdBCRGb7UKUPyk44FDkT2YDmeDEQkAyIPTxFl9fXl9swtypD0GsQuBQ2M5aTiILMYSDQ
5pKQPQn9H3r5FRhzQsaVnCQMnLBI5lB03/xnWqmIQ3+1ljaidvFlsODkTkqIryvzzPaoLUihWvAv
lV1lPsowNMqJgcut/Li80P54BwYtQT304zxJDxdDiDQGOO5a54b7DqqLnZKT+fL7xJJAvC8q5MHl
3+rJKpwWrSDLq84icQI8pk3yjWQ3bVoC2dhnZ2wyyyO9BJo0RmtitdkavtK28LrGEQfdiScFJaHv
AjpoAnPpXOdl2nNSy56aA+GKfvgOW4AgydEKXwqE3Sw2KR9oHtLn5ADYum2yS8/AX4j62Nl/iIwL
2DfHIB4/kivUVKRmj0ADjqojrTLKLXCEn/yTVwBxV7kfQClMw+RRZGZuTlrpSyiu/GeuLuLGo/TI
w5hm0fAq3qSbpkK3ZkALCdTPrJEMi5Ye6yrIn4Cl/RK9Olsn5fr7lIBo8cugRjeedQW9V0QJrAAV
vXTXRWXRnm8hZ3W/NC8TgmlT+6A4qUp1hEwHItigGEeJlnt8o482DjXstcPX5/i+Jmy2lPfW2ueT
rH1/xJIBqbT1JgQdoiiMXJiksW3qdvhnaNuVkdQP7OY+vf2sE2KY4rO4oRuV2PJ6yFyrp5o7vNmo
mNl8xHC+mQnvbmhiSjNtTJ4O30JI7zEVaKGzVlf6eGowBjaffc4ceewz8EL2vhOmzyYgcyZa9hS7
jRsiKTwFXi8lGMKL5Ju5x51TOhGMWVEvWBoy5Ampi3Kw7PgFwJ3Odb2oDP+MlynntpEE4P9wJycc
Q7ZnlkK6Q0ZQYqV+DMDx77hg0CVbM/c5yutOH+XwasBLu5mt0hF1mkIPryaReyNmK/kEpg2H3zJz
wEtQEJBAcQ2xOhK0uQKQ5HZipeBrSnu9pcrwjI53147dVmoddUfWheHh1uf4WDExXFXS6hFlQwbd
nKrY4npPeMxzit8lFmHoJThhdK3yE1pFekxjr/XwjPGcuo1cQg6cNXMudiCSFIpSneTfRfdWmgYN
9UrhRprriGJlnETpgg3TqWCOPzw/CN/QEIdQwUdZVm9fjen6iaAuTHhxjnnTs7mIuFNSQ4W1rIFC
eYIrklDLxnSiIYI4nvczKajth+FObvXZ3n4rYDeLzCt5cHNf0FHeTqzVtthrqc92nNiwhaiUoPkV
+iFy2uR7niMmqBsgk/xl2U3bG1J0nFIf1XDHhRugxf7mrpJN9fr3gZgbePQjyET3qAlcFcbxcsDF
7A+ROkd3XYPj35KHV5HoZCfHcFp2rvllZKctSF32mEndD56Aw3ygkL8+XaUNcbXfj1hJGNpFtMlF
VgGWtzPVcj2RYitRTH8qpAnfFw4S7W4FeiwFohc/ROy0kntq/RUHQQ/xEDv1tDmQ5EhafxLAdJwl
J960hC3NM+GmUpWuVwuMVN9GipPXGGVU/F1E4kpjFT39Fju1Lb+1dkoENv5KEneKChk1Y5ZFpAbi
ztsnffSbSseimm2RJr10zpzi9w8aQd7cCfLkrOMxwbClFi9mkljZTN9H+QQ3fhXg99OmnmXRxmrN
DPAH7pFa9HIGZB738jZ+0OCTpSn/WWo62U7Q4gC+DVoLIvmvkPAMQdvU1BBKquVMApmHg/7e5aww
txj0KusImrpcPzJlCwKRnWuGEJAS3B5DR+L/IMuhstNaeaopYoBHAaI0FQyDiLUj4Tr9Wp/kWnK9
WhdIvt6BRCfsGZTY7AVmuZ7d9FL4tZIJeUnq0I4V14aL/uRLetXB0hBsQYkDkgIqI4F1bz/yJSvI
uBkGxxTGUymT6vU4fuDB9m8d1JtrsVr7VqlsGTXi+UrFl1hx71eugadN6WthTttgu2oJDxL5BMbb
XONx9CQLIX7fS/lFo1qo4nkSuBe/I2r/2oL3s/zKccGMa5YR6GmyA68vEdVyj/5hDz2eE8zXpvIj
QBuMItMuIfJAeuAktZG+4cbj9g1zWiQT6PLNU8radALP0Wr3KRqZNPg0mrgcpDt70GJ3HxqUKsFi
GSO8tZ+rDg2vWm1dKRuwbCeDfNRMrvkC7/3YhcjUjlzqVqjjB4BuioGo/685a+bYLxbhVzPMNlfJ
WE5nL8tP+CWmztAzVu3C1K5+WQH/Qd4IP3IdCwW/5ebvJjyzskQ5gozC4lV9U9Dk34dmvHsyZF5B
2ehNAfyBrjt7FoEJY3q2B8g9kudHJ0bCasSFHZYdlzfuPaWbd4ABQFCc3wIfqxE3ATbbCTO0LLeo
SSxKtwxACow0osnAzCnPp/TsOIdRP7Ph8Oha5eDkMkt7VYpRZxBDWSnRHKkKRXMXvTw2lH8qprHW
R2z82PYWqFiGm/HjxmDzfcrc2MRyCYktWbJGX5V8ObveTMd71/N0vJNYHvvwkLRbgBxEM6O8fI9m
HfewMxbgo62OLUCUWuaRHm1K7qZfi6Mx8OfkI8TE9ZKeF1M48fnHQC0BhLRy7UGhXkHp8E5qJCab
3sp7yF2FFSmrgpkWaIeArM4SM+yGp68EP7AtIqMbYWiGlE9DqW1wEwwm01ECMT8hWy7iTzLHWW5K
SNS/NfsqLMIVOHp8kZH5Lz2AYydpF35+9hGFrSyuLmevgtMUMVjUTw27fqPZ2xn/xcL5NLT3Wikp
4vz6GijlGu5W+8GrjbYt4XFP9SN0wyO94iDtBISRHvXaBa4au54ObY5i2MwNxnUpB8D9DvXXj9O3
JN6F0a0/t5cnn/KJotogdiaYHvGC1n2+iB8VuLkK3JJ1+mAryxk8FBc6oNoXTX0PbusbnFE9bcr6
gfj38LLPWwTGZxNuSpCeNYmrOkH2rl9qVNpPhpEORYonUHPIFfwf7H2wAqmMrKM4XES6vo2N/3mf
awjwamIMrWNdfUxfNgi555Dq4u4lnC/F9J7kD9GrJi2BDjNsNgCpsUTAIu4vadgDts/K/MRKa0jt
ky4qHZND7gZhdFJm1CuS9zdZ6VZxWIP9cISoOVtz3xK55F8ryh7Mqu/sDNU/BZ/AUbFTfbdjsBnf
Z1HBhQ/E6/g49Qh7evFs+JjeJbrD6sVqaSS+80dHtzIqFAKQdPMr7u5O3x4XQD6wPJhQd5M7YRBi
JmBj5zrhKLeqanNuGYvr1sYbWLulN9dpOHi5+eyHWYke4wN3LjtXcTvh41QUGtIOF0LeBrzj6Xz6
kqsFhR69VyOGICHZM9Fd0LDvo78qPeDmxISNNVXXB3V926A/pIxXd1JE7l7F59DfGGx/YezaW1Wr
SDU8BZ6gq7kyYzFMHnMqj9kt7LNT3vEng4rqU0Y+JL6F67EGXKvf+jfM2YAIpNpF3YCKUAnsn1O3
kkFnEcotjw4QIHoIMPmrp7tAtY5AIUVYWfcWtzjyJNfYSEhky06GYy3RkoCif9CPiT/DqV98fTsl
uIGuQ0aKoaUolKxCzTeIucWGKtAspF+mT4bEEnzWiWh0MZ3w/mcV/enE+H9tPeuiXtvocZFI/ox2
aegKRfPZO63jPplNGfYB+qRIzVLUjVHCEukZZRgVaIUjHOmT1jfpEs/8QINeNq0t1IyLwClAf6EB
yJDeNky00cf93cat5KW4eBXwu5lle8Vlvf0Y/HnfasaslMC8WU7f1ycpYxOiR8IBJQ7T4qdYO/YF
zHPftbz3whC3sF/ubbMfNazcxf3X1b3ZAZGJJfxI6cPxMNyLbAfD0scizGh1JZUAqJAVXPsMT/Mi
rcyvy97TUw/tO2tUAqMwW/NZY/xGJgAuqJ2M37Zf99TIf0rb1RGQgSQKxXV/npRaThq2ezgLBIuD
ZAotNuS1en5BMcpZE6cmDtZKY298LizC27n/qXv44JbQZaajoeN+91dy9eHANIQHjui7mkMGbn7q
HNRgJVcBjKgNzGNnyUDFVSF0PXiGz3lQtXXeW2knReiq0kQD9qPrHrz3qP0os5PU7p/7CIsDBhGT
hQJfUNeTwT/JJseBZK8CJinF956dYqvolq9jVKXOUPu4oY/mMt3NaQJpqQ0Mj7sCP4u10ymaJZBS
K5suwglLcKJkXVHxVfsEwV+QrjqttwJzThOhciJHdaCczG6P6dLWb1mKDxD58cS5cqe11fkcwSuO
PzGiGcGd7Spq1Xsz0wJQ+6UKo85JesQvr8ZuxdF85Rh7Ll2oBDIi2OUX8Ak71qw9R+gYT0uagQip
RIMQl0le9CE6a60ojMaXv6bCiz4AdDPDwe6Wv36ikRJ+E7PHs8NpnJleJyFJUaIjTUqtWidv7F+K
Oxwltx/k6oaPUBGrY1aQLeEH1S6S+gdR/kYAvsyeG7Ls++Kv9sN74mWSDAvG8AhuNfHdngkIG5tX
vqQvmq05HAYVeBZzT9FnyZtaYc/1l6GQXElr09+0sX2GwkNkkr08YbixNd30ei1+SpO+nCEXFZ0U
0a3yHUxhMBAeNrrYRg1wSNcveTzPBLHZmoqOiyP2LC/a7oMWiSYmLSE9m7O3x6nbAcvddkhftWIb
3nC7MLrvXWJifCYhqkg2LPufs6Cpv4i1TCvy+aoxI1SiVeanyjslcIZzYNcfWeVS8r+maeYmC0i+
xaIycHdsCBzck+BufJFHhhTP7RQp6xeZq6Orrd+6goXjUs5sNu/u/mCJJ6T+EsdfS6U6qFwlN9KQ
JGjpN9ucxsydvgzOWDb5f1w7xX9LtIW0MDTZEBzZzlMlwbjMTv4I4Mt1RP56veAAKjVN6vZ/Odom
88/7OFTgBwlGcakrGucZ6sElhcg24fXJVYZ8P/fh42dK4IGDBgj2NqQRMhXFatggAjxFsbn8ymsx
UrawCyRw2JD4oqO1gP4ws9hyUIWrm983q96vmFagbjS4wDTSEb8zVki6oeLqmpmIEuJ0ciEApLiJ
lUpCn4ZseJ5/wpeqAgRu08+i+FWDu+Pu7KfpseCWLorF+PyUZ1goRaQVM3pMKEMQnnRmksNZH9C/
Pul1yVLxYQvIOj6FPAxxHiIvu+Oa4pfTBBVdF0iQzG0QVljfVd9eE/rBjOyJhhw5lNTGL6RSIcQC
WqCGhJkYo7XRl/Zt+UTlPAdpMOa03csX5OlT7Kl2l7I6lGhlJbW0vOAUGD+dHxi3Rv++pFjb4Xnl
VJhzizRkIhqSe6e1sa5OiziUdtvECo+hWn/jiZoc1dVJ8C6kIJHPWxLVl/tbxQuWltpnsXqYYWpc
vRbRz+5ILmE/UacBSKeeuxP/iunfCodV7w5Q1uy/uMKYpkPLjJdztlMGrt20BA3IYDqAylOcssJZ
A0/8+9lhdJkTeLBtTlsIXaSxh1qiy72ovnu4qrHnaeeoneFgAS1jXRNFLP1tU24PKUE5VGVjZF/a
Ujh9qbwVrLBeoops7QEER6y244wDQoWnHWk8ejmsE2l1cFAShB3xDuB/+tmkuthjK7lHIN0ieqkd
0cwa7EK6N319SgAOuctu3PnzAcK43PxhzQ76mn1vsTZkxGFdK8bsfaOUJAFw4rAxQ5w+X4C0Zs6V
DNFXDsZ5Wa+R8SNRrF47U3/YJnYfv32nGm/H7ezoHKDcH9WeDe6F0hZbl8tanFl3LxOBRceFpmMY
JMtLZiqjBst3dLECsYx3Gimil630IvWZfkdFCNlWStjEssAe1rqLvLaoEKtVIDM1FDxWMFVAGNYQ
vl933ZcUF5H/MX6GxdW970u18OFTKdNnWjr50wvujqo45HER1B5dzDR4R7UB2afxZYrzjgFRHuNa
s5DQijTjr9nh6EpFt/0N8U/zpeERHAKuL6sKT5QvjSzbNKziluRA/5DOmV5Bc4jq3DXZlxj9HYer
HjyXN3UV2M276uI/vUpED9ckkrZk4GVCgyudqf9cFA0f60X8K3zWDUlNT0AzbQYcqxL7FUify5RC
OKhv5iDDwJOTrfOS4K6Ik0RSen8C4QejqXNH6Z3ERt4uLt/SPiBTskoeXkxzhc7NL8btgMIHsbPr
Qm+nwQXEd8ofx0aiO3s1qA8b/ZgMl6jT2tfBRbRDgpM1CFZJNxWJV9Lh3CvIEIDeNCbNnPPSaEdK
3OLC0Lb94He54HWOK/U2h5YEro0a9uA3iSjXvXhAzivM8l3N6JHlPI5WWO/FwZslps5Kb6cdLk/D
/sonAbtfjbGgVxlQSKTD7boKZ7UVDaympRJr3QA56S/xwc34v7b5lmFcC85BUHk2OZ8XWXtQzBBo
x2Q8iyHAS6InymXhCCYIpbdor59YSVu5SiALaNMyGx5scyCrs0pV2yVaq+Xei6Bup0FNipFFmu1k
tXpjD332npQ3v8SxdP7tAL6Zl9y8gGAbzn1e3UIvH0Ki4pHfV9cyN9NzCe6Il4W2RllYwlmhZ68n
mk7NtQhn6eCQNy7pEC2c57VmojNGwnCJdiUt/MrAXT4jz28mZyjVZVZ4Fx+9JsPXu6yynCsSHUvS
zZqdmSwe7Ru9+3nwriG6tjT6nhmC7ZBLHPGBoGH75IbJ5FiBXB9kvWC4JMt3UEwdaXo3q1zoeduB
QgG0EL3PEKP//9CgkMrW6Mcp2bTEeruyVoe/5rRuxeaFHUeDHGJUlqbWKV71qfiyTDpicjNkOPGk
1R+bPF5EXn63+CCiWEHWlkJ7PomqIMdbxO85sAGdkCDSicQqC507gBMqhafsZ6rwH+obc4pQPPB8
f/n2fefMW6OvqfKpcLk2J2EjbMM/G5GSkuPoi91CL1zRMtc4rdRrx2IxBkYZG52tZL+DX/ffw25/
cJ5uHEV+mlOV5Td9SPNXX/dK66cMLoxASvhq5ekj96UbB5ViuMqxqOYxbnasb9MhowAy01yXo3xd
AbLYBrnxwLtIPw1Ch1u2Ttow5V6J0CJ6gL3tDhIvKbOENHN5A5dK7QfXtdbiuZPNr1nrj8jtmDo+
uHOoXN/F1WluJQ+qMQUaK4HHNuc3g9mDG1Ahd4ls3djzdZL8t4GwZkbEdoJ+gAFeWhAQA/5mjFYm
7jbHXWpPplnX3VrI9+MP/w144ymTYKfzp/19RWXlI/Wl5h1iHxWKIW657N6U2aypkQDdgCe4+nbn
IcRvfu5OSbwN2lJbL+wu1AHcdaIm6D/qoY8bT/zCbeO0HqXvdO2p14g0nvdSG25TBrA+76JHGZ3A
TuKHF6yZfuTZQFwPMoR8sy2FPzNQRl/EQ5/+cBzhoSqPa49deH7/caJ737MnwdR/Ut82io04eAWK
5sL5P2mYLiLz2K6ciJ+h2m7voGFnec+qyFSH7kJ9eoei03dyjRgVpK/Nek2f3xLAvqvV8UJXBgKq
H2hywu0AHoXS3yhb2c6Zgv/V0A0rmcCppLGKDIz52B08Mnp529y/tM8ifhWxeo55KQYI12CHoHSV
vwR8rI9l17LNGHME8rgqEro+FOYzVtMrQpz0t3T+JIoPCgdpmdITnfU/gjo45TNJnP/jf9IYJTQL
fbQp/PVAzf/FqjAbb+kfQNvCbOwQNdodTa/lP3ZMtlPeiAlEJ5Pxsh3TcIa+Gm+Ad/ckhmCKq0HY
Q1VR27efNSPnMbMuAj3jPyOHmflZ1YLOiPMW/iW5k/DybkqENnM68Vx697/I/xDpV2W2QJFKmNz1
F/kAqDUMlE+dxAqY2mXVeZYKWzHz0ik1YLf8a66ciICUTinNsdtegzN++tAyLlSsSlJQWwcCWMGE
uYsICCPRDYTnxz4MBB32AF/GLwpUnfVQmRXPr8O26tlaP+/xlJp0R8t6HH8pqJRxhlKpUE54V81R
z5GXIOslixSXe8GBwfE+hx2+FpxthgoEZxYEUuHSnp3iiU8g2C5SMixuG8lupqtlfaK21kOJ3cXI
bUIVfqKmz1oiYqzC/4l16L3VestLopq5KcRY/jaoLaFvMH9ML917LXhOc98uXB6EVuvJ5c0cm6jW
q8DrpMJ/2/9cPpWzIYf6w8ZKYCbrYWAk7N8lhs2OyDI/Owm9Z8XktuolEeKxWQ64tXwncyAGqiRz
axCAPyFN/haeD3sOoXciozFbG7cjs4shHG4iSSEl0QQP+OYKDAhmUWd1fryftiiFAk2Ao3xRLO1F
ezI1eB2r3G0lWRvoKi/HbACxbulE806UYuLPucs2F9QBFgWqWfI2tpcGKSOk1Yygt0psPeuh7Sfn
3uYSbRl0DAq+xsk5dFOmKyW59kx4Db0+sMvI52zM0boKfKbkRn905/pVpFmYMoiq/D0dFpgF3cXb
SKbu+KDqi/qqSIP3rNI9DIZHF2B9F3rUbnbEq6h08+3GhtO3nNU6DqKgbXpRxNxcK0xxo1mETxCa
LCa+6Gye/uI19KzadA6ACuqZyCBfDHoJ3usGSIw6brgLbAMLPmjgZEVYFA/xCEMfZQ9GG4wOnRxo
N7cfDe/Tz9WTfvpUszTDH4/5w0fF7yZoHr2tGbqOy6zmdQFC2hBOSBR3W2pAMKBE6FJRS0+rVszt
uYBvY1BeqOjbKx+O5cVxrHWgG8MtZAMeK+Y7py35kg+JH1Lx8m54pYJBQXe4rw555ZgaTYM6366W
FNT899hkOyH3DRjhr8xVLUCBwi/oz7N4/oQVh7DGisWDp+gm3Q9R1MFtCtwhrJSEODsuv5p2kl18
mij2dXvCYumgGoEMlJ5cYdvVAziSqE9blQ62M4fHITN4TA89bllJbFnOwVV6bA+3EQql4eKESyZD
eL6+URdYlnRv9HQX4M6EW7gJbOOQVV3v5dpX3PX8O+zpjPyGR7e6iFqOqZqRnegs3WBmsr7TIG1j
vj2UBNv94ys46lnGhCVs73pY1OudscmLWphJCa+8J2xk+JCGArpkfH84p1ZCvKdLgHkpep1bc+Be
EpcaQgX3oVxKXROJB1ddfp4dnMoB5bPMxcVatWyU4muoTIajl5lte+GOu5BKXw65bN+OQF1bLIej
az0Ziw/t96PinaL9r0LXy9OlAkdWXBpehGbnOUT9x4TY9cG2sbUMhu5fH2tmddLBxdDlHUVPVLGQ
NQLMejJf4XU+pRATAXOuy22t7DhMD8rYdyDZctSYZtfTDiXbAQE167E/56+DpmEorf+6Pc/gHKhK
CycMIdvdlokwbXJsyqhtT6G8HO5JSAtzRcXR880VOz6poLoLu8E20KjM2tf4Gj7TXiHGac0AIb8g
V87LU3t3l0rfzA2XWYa9rFxzecjEODMkYTYsdqEJi75Su+nSWBMEGZwaN9NpjRy7nsOGxc+rqviq
V4Ma+ueGCw0bwtZSpnDZt6n+D28Gk/dKqgV2pwaXTnbaSiNS3Cm6kuIos5DvmVcwXww+33YcCuWV
wmFmu5ZZ7JXYH8pnV7Jl6m7iaxn08GgOULodOyfvSv6RZ7zHghcaxv9n2Hmb8FBtZJn8qbNW9J1U
014zhO42Upn4J9RtYgxpOjsFHFvDoxueLT3x43tUq98xleCMD5gnlzaJgQDPPCKhm7B9Kz/473rs
0ZcIH08XtfQ57khP2sb7K5tqTojSSwhI23ofbjiJD6DBkRfbvp5/AD48zjqP7kqE0bTSao9/EqTN
JWi8F8IjYRXpXwX3/GNIU3jIly9XloW+Sw6QjDE72ktfFNiIWFQLFQ6Fjm72eKVc4mSrDv9PBJbr
TZKSync/qgYWbcMea3hybKORcb/tPJ2FaqIja8tS1PvrNxmhVKx3j8nMTN4LkilMQNobkflW4Eb0
oMmn6P1rq2Q31TVGoy7zaZA00ob/t1CLSWxeep67EepymVKOWZ8ZcXdDRTUc4USe0NifktNNiU4X
5GYeMbB4i9X0yRoNzIuA924mZPP5z8geBmP+foWlXKmiIzJoZtJPCdi1HA81xOOd0um4j7o1Dobd
mMoC6112xbLT2LaCZeUqWTZmx5/WjrjMG465QWU2ySvn8Yp3FrM/IA3CQNDyvYQg/Flxgf0eM36l
rqau/BqIKyRwVh1dF7p4Yvr09vf39EerE9sNbI8KEygq4c1HQ4Xe53nmhalwAlaEjv9c1R/Rt7sD
LasLvUFHqw6cBv37+WmS+z9MD77Snp/B7dwQEX3Jv7ZrgYnYHr8R3+VY+aeIWgq7FMF2m2scfDJ/
XUarJnM0eO48ZA8Q21f0Hl+Q7J7ZAoSzSVCPKOFNez/zWII40RtfZPqquQElrfolbGFH/nxEJbGj
5QMnxsz1G+swetdqDEyssCn0JEXRr5Miy5CRhuLPdk/HgdMWG8YmSE3uLR4/kZrvFuQ1VTtsRtVQ
CUzcXWTElVUNTRFNnMb1SoE6EhfJLVvXMVyVH0O4aeE8gqFoBvdpt5qzhw1iAeujnDMMOLphEtw8
FDqKgmSsW9uX+ewPlPe2BkLHsO2QE0p85O74rIItFBjed4j79XWI5bAVn8SiZuk8KR5M49gHjUHz
IUlT0Rhv7J7yFxU/wojIQV5ql1EAYcpT+R+xB6LjxQnvm9rKiumXj3nfY8JMmBrp/HudQFuRK4gf
T9Q1JN//EBjEpE81+7/xB6DLUY5nWTea0BStcexmJkQzyaamlhCOtETXdDuzOg7oNQyuPfrJz2Gt
VOBotmY3MxjbY4PQro/dc9yHaYsyYi7tdpc/v9fIngniwoKucZvWJInjWjUt0a3uWcZelcweysvb
7FIsYEvHC3bnU03vVA91onOa6+i0aI5XwUvVwHF1LPFQW0qVkLUnY71DWRVPapc0hnlwAlOSiSV5
Cq8/nEkZrzGpeVd87WzHr7VA/fTj85KDM+tGhKyo73O4q5uw9iXpKzhZkzVO2EMPH3N6ikqA12mA
3hj4DJOc1DqmbG3NVFGjA0Vl3vHRNCpD51wYn8ED6lHy09PfYsXj/Bj/m7PGjzG1ufxb1CX8a38x
H9w36DsjpxNqUqRhrKs6uKS51aPdfqbgAiR0MpVv3GPwIrJInoVQdxZAEF+eZG14xt0EF9K9LhXu
fLzPmHoLoaUIl3gaKQY0o/aCi2n3rImLNcF4GUXAdiNgA+FEE5eIX2cnNE+7uKky0NhmzIBE+wjj
Dj54xCA9PocxFaohhC8iQ7JIB84VYyYlmeGCty0Zkl5QB/awTjE24F+FjCux8Z0APjvgwCyib6FJ
PW5fBuOz/1KwqmvbZxd0MjFXPx9QUYogdkemltEXQMIsVzyYjucXXgyaowCNG8QTDxANBu5Gmio9
j5iZi56/55EHVdONXbEuYqgkjgwii7okT3+uwFz7QLRVW6n5mEAacy/mM6J1/xaGXZg8g/FtBkkG
g6he0xAb2fnEK6QWz0NPuHGpfv/+Aov6kDiIgeHRwXJRdt/zMC8GPQhMdv6XuI0akX21H88Sw4UU
DypxCEt/ODSsnIlCpLIDT9b0GYFTm9YRkZ0rIOi3lSR8u1jQ8mHWyYv7KMJf4y0zQcc1nzzQGYcG
vlG1B5EYJZ7UzUUMLT/AZvGClBwsesLXDIp8MzeLY9v5WjQun2kzfHMcVigLIrHNNeq64C8nZHLS
ELowM9IwbQ58E70SA7O8SNB+LBcz54rTa8IiAP9q3hC17rsFGwl2x8pOD1ytpjJw1bHdT7pZneeR
GgFukkXtB0aukl7gadrRxqmkbQqIuHeMZJifFWIVF+bktmVekoPTzivHWKXZLT76QusrZUeMyfko
j6LZoLfFucUC58bEEE9SVRv5s/wuZmZihbAx7QmTWHKOXfCIuQ1xNTriQIhUWCClnF6gQXB76w7y
FJrSi8gyWT+a0Nzfoixt7kYQvdiE7ZmhIrb6FxM3+S7l2P8LtO5y/tgQ20xWQ537o8GMhkg8c8rK
eockwjqV9IjRdKMFYvIKcKRKtmsLaPNniFgzqDJNjftcdk/LMM0jQvYwfqK/88IXiPaBIRT8NH9y
mojqAYdDejpt6GCoa3U/KjOKj0scIPWVFv2BUUmSAsdKT8LC8t7kOjfgyE/5nbprZe0Nu2Yzb4yx
a/wvoDgXfINeef7Ms23iZA/EGxBOIlD6K7zHcAC0e5AReT1O/Q==
`protect end_protected
